module AddRawFN(
  input         io_subOp,
  input         io_a_isNaN,
  input         io_a_isInf,
  input         io_a_isZero,
  input         io_a_sign,
  input  [6:0]  io_a_sExp,
  input  [11:0] io_a_sig,
  input         io_b_isNaN,
  input         io_b_isInf,
  input         io_b_isZero,
  input         io_b_sign,
  input  [6:0]  io_b_sExp,
  input  [11:0] io_b_sig,
  output        io_invalidExc,
  output        io_rawOut_isNaN,
  output        io_rawOut_isInf,
  output        io_rawOut_isZero,
  output        io_rawOut_sign,
  output [6:0]  io_rawOut_sExp,
  output [13:0] io_rawOut_sig
);
  wire  effSignB = io_b_sign ^ io_subOp; // @[AddRecFN.scala 60:30]
  wire  eqSigns = io_a_sign == effSignB; // @[AddRecFN.scala 61:29]
  wire [6:0] sDiffExps = $signed(io_a_sExp) - $signed(io_b_sExp); // @[AddRecFN.scala 63:31]
  wire  _modNatAlignDist_T = $signed(sDiffExps) < 7'sh0; // @[AddRecFN.scala 64:41]
  wire [6:0] _modNatAlignDist_T_3 = $signed(io_b_sExp) - $signed(io_a_sExp); // @[AddRecFN.scala 64:58]
  wire [6:0] _modNatAlignDist_T_4 = $signed(sDiffExps) < 7'sh0 ? $signed(_modNatAlignDist_T_3) : $signed(sDiffExps); // @[AddRecFN.scala 64:30]
  wire [3:0] modNatAlignDist = _modNatAlignDist_T_4[3:0]; // @[AddRecFN.scala 64:81]
  wire [2:0] _isMaxAlign_T = sDiffExps[6:4]; // @[AddRecFN.scala 66:19]
  wire  _isMaxAlign_T_6 = $signed(_isMaxAlign_T) != -3'sh1 | sDiffExps[3:0] == 4'h0; // @[AddRecFN.scala 67:51]
  wire  isMaxAlign = $signed(_isMaxAlign_T) != 3'sh0 & _isMaxAlign_T_6; // @[AddRecFN.scala 66:45]
  wire [3:0] alignDist = isMaxAlign ? 4'hf : modNatAlignDist; // @[AddRecFN.scala 68:24]
  wire  _closeSubMags_T = ~eqSigns; // @[AddRecFN.scala 69:24]
  wire  closeSubMags = ~eqSigns & ~isMaxAlign & modNatAlignDist <= 4'h1; // @[AddRecFN.scala 69:48]
  wire  _close_alignedSigA_T = 7'sh0 <= $signed(sDiffExps); // @[AddRecFN.scala 73:18]
  wire [13:0] _close_alignedSigA_T_3 = {io_a_sig, 2'h0}; // @[AddRecFN.scala 73:58]
  wire [13:0] _close_alignedSigA_T_4 = 7'sh0 <= $signed(sDiffExps) & sDiffExps[0] ? _close_alignedSigA_T_3 : 14'h0; // @[AddRecFN.scala 73:12]
  wire [12:0] _close_alignedSigA_T_9 = {io_a_sig, 1'h0}; // @[AddRecFN.scala 74:58]
  wire [12:0] _close_alignedSigA_T_10 = _close_alignedSigA_T & ~sDiffExps[0] ? _close_alignedSigA_T_9 : 13'h0; // @[AddRecFN.scala 74:12]
  wire [13:0] _GEN_0 = {{1'd0}, _close_alignedSigA_T_10}; // @[AddRecFN.scala 73:68]
  wire [13:0] _close_alignedSigA_T_11 = _close_alignedSigA_T_4 | _GEN_0; // @[AddRecFN.scala 73:68]
  wire [11:0] _close_alignedSigA_T_13 = _modNatAlignDist_T ? io_a_sig : 12'h0; // @[AddRecFN.scala 75:12]
  wire [13:0] _GEN_1 = {{2'd0}, _close_alignedSigA_T_13}; // @[AddRecFN.scala 74:68]
  wire [13:0] _close_sSigSum_T = _close_alignedSigA_T_11 | _GEN_1; // @[AddRecFN.scala 76:43]
  wire [12:0] _close_sSigSum_T_2 = {io_b_sig, 1'h0}; // @[AddRecFN.scala 76:66]
  wire [13:0] _GEN_2 = {{1{_close_sSigSum_T_2[12]}},_close_sSigSum_T_2}; // @[AddRecFN.scala 76:50]
  wire [13:0] close_sSigSum = $signed(_close_sSigSum_T) - $signed(_GEN_2); // @[AddRecFN.scala 76:50]
  wire  _close_sigSum_T = $signed(close_sSigSum) < 14'sh0; // @[AddRecFN.scala 77:42]
  wire [13:0] _close_sigSum_T_3 = 14'sh0 - $signed(close_sSigSum); // @[AddRecFN.scala 77:49]
  wire [13:0] _close_sigSum_T_4 = $signed(close_sSigSum) < 14'sh0 ? $signed(_close_sigSum_T_3) : $signed(close_sSigSum); // @[AddRecFN.scala 77:27]
  wire [12:0] close_sigSum = _close_sigSum_T_4[12:0]; // @[AddRecFN.scala 77:79]
  wire [13:0] close_adjustedSigSum = {close_sigSum, 1'h0}; // @[AddRecFN.scala 78:44]
  wire  close_reduced2SigSum_reducedVec_0 = |close_adjustedSigSum[1:0]; // @[primitives.scala 104:54]
  wire  close_reduced2SigSum_reducedVec_1 = |close_adjustedSigSum[3:2]; // @[primitives.scala 104:54]
  wire  close_reduced2SigSum_reducedVec_2 = |close_adjustedSigSum[5:4]; // @[primitives.scala 104:54]
  wire  close_reduced2SigSum_reducedVec_3 = |close_adjustedSigSum[7:6]; // @[primitives.scala 104:54]
  wire  close_reduced2SigSum_reducedVec_4 = |close_adjustedSigSum[9:8]; // @[primitives.scala 104:54]
  wire  close_reduced2SigSum_reducedVec_5 = |close_adjustedSigSum[11:10]; // @[primitives.scala 104:54]
  wire  close_reduced2SigSum_reducedVec_6 = |close_adjustedSigSum[13:12]; // @[primitives.scala 107:57]
  wire [6:0] close_reduced2SigSum = {close_reduced2SigSum_reducedVec_6,close_reduced2SigSum_reducedVec_5,
    close_reduced2SigSum_reducedVec_4,close_reduced2SigSum_reducedVec_3,close_reduced2SigSum_reducedVec_2,
    close_reduced2SigSum_reducedVec_1,close_reduced2SigSum_reducedVec_0}; // @[primitives.scala 108:20]
  wire [2:0] _close_normDistReduced2_T_7 = close_reduced2SigSum[1] ? 3'h5 : 3'h6; // @[Mux.scala 47:70]
  wire [2:0] _close_normDistReduced2_T_8 = close_reduced2SigSum[2] ? 3'h4 : _close_normDistReduced2_T_7; // @[Mux.scala 47:70]
  wire [2:0] _close_normDistReduced2_T_9 = close_reduced2SigSum[3] ? 3'h3 : _close_normDistReduced2_T_8; // @[Mux.scala 47:70]
  wire [2:0] _close_normDistReduced2_T_10 = close_reduced2SigSum[4] ? 3'h2 : _close_normDistReduced2_T_9; // @[Mux.scala 47:70]
  wire [2:0] _close_normDistReduced2_T_11 = close_reduced2SigSum[5] ? 3'h1 : _close_normDistReduced2_T_10; // @[Mux.scala 47:70]
  wire [2:0] close_normDistReduced2 = close_reduced2SigSum[6] ? 3'h0 : _close_normDistReduced2_T_11; // @[Mux.scala 47:70]
  wire [3:0] close_nearNormDist = {close_normDistReduced2, 1'h0}; // @[AddRecFN.scala 81:53]
  wire [27:0] _GEN_7 = {{15'd0}, close_sigSum}; // @[AddRecFN.scala 82:38]
  wire [27:0] _close_sigOut_T = _GEN_7 << close_nearNormDist; // @[AddRecFN.scala 82:38]
  wire [28:0] _close_sigOut_T_1 = {_close_sigOut_T, 1'h0}; // @[AddRecFN.scala 82:59]
  wire [13:0] close_sigOut = _close_sigOut_T_1[13:0]; // @[AddRecFN.scala 82:63]
  wire  close_totalCancellation = ~(|close_sigOut[13:12]); // @[AddRecFN.scala 83:35]
  wire  close_notTotalCancellation_signOut = io_a_sign ^ _close_sigSum_T; // @[AddRecFN.scala 84:56]
  wire  far_signOut = _modNatAlignDist_T ? effSignB : io_a_sign; // @[AddRecFN.scala 87:26]
  wire [11:0] _far_sigLarger_T_1 = _modNatAlignDist_T ? io_b_sig : io_a_sig; // @[AddRecFN.scala 88:29]
  wire [10:0] far_sigLarger = _far_sigLarger_T_1[10:0]; // @[AddRecFN.scala 88:66]
  wire [11:0] _far_sigSmaller_T_1 = _modNatAlignDist_T ? io_a_sig : io_b_sig; // @[AddRecFN.scala 89:29]
  wire [10:0] far_sigSmaller = _far_sigSmaller_T_1[10:0]; // @[AddRecFN.scala 89:66]
  wire [15:0] _far_mainAlignedSigSmaller_T = {far_sigSmaller, 5'h0}; // @[AddRecFN.scala 90:52]
  wire [15:0] far_mainAlignedSigSmaller = _far_mainAlignedSigSmaller_T >> alignDist; // @[AddRecFN.scala 90:56]
  wire [12:0] _far_reduced4SigSmaller_T = {far_sigSmaller, 2'h0}; // @[AddRecFN.scala 91:60]
  wire  far_reduced4SigSmaller_reducedVec_0 = |_far_reduced4SigSmaller_T[3:0]; // @[primitives.scala 121:54]
  wire  far_reduced4SigSmaller_reducedVec_1 = |_far_reduced4SigSmaller_T[7:4]; // @[primitives.scala 121:54]
  wire  far_reduced4SigSmaller_reducedVec_2 = |_far_reduced4SigSmaller_T[11:8]; // @[primitives.scala 121:54]
  wire  far_reduced4SigSmaller_reducedVec_3 = |_far_reduced4SigSmaller_T[12]; // @[primitives.scala 124:57]
  wire [3:0] far_reduced4SigSmaller = {far_reduced4SigSmaller_reducedVec_3,far_reduced4SigSmaller_reducedVec_2,
    far_reduced4SigSmaller_reducedVec_1,far_reduced4SigSmaller_reducedVec_0}; // @[primitives.scala 125:20]
  wire [4:0] far_roundExtraMask_shift = 5'sh10 >>> alignDist[3:2]; // @[primitives.scala 77:58]
  wire [3:0] far_roundExtraMask = {far_roundExtraMask_shift[0],far_roundExtraMask_shift[1],far_roundExtraMask_shift[2],
    far_roundExtraMask_shift[3]}; // @[Cat.scala 33:92]
  wire [3:0] _far_alignedSigSmaller_T_3 = far_reduced4SigSmaller & far_roundExtraMask; // @[AddRecFN.scala 95:76]
  wire  _far_alignedSigSmaller_T_5 = |far_mainAlignedSigSmaller[2:0] | |_far_alignedSigSmaller_T_3; // @[AddRecFN.scala 95:49]
  wire [13:0] far_alignedSigSmaller = {far_mainAlignedSigSmaller[15:3],_far_alignedSigSmaller_T_5}; // @[Cat.scala 33:92]
  wire [13:0] _far_negAlignedSigSmaller_T = ~far_alignedSigSmaller; // @[AddRecFN.scala 97:62]
  wire [14:0] _far_negAlignedSigSmaller_T_1 = {1'h1,_far_negAlignedSigSmaller_T}; // @[Cat.scala 33:92]
  wire [14:0] far_negAlignedSigSmaller = _closeSubMags_T ? _far_negAlignedSigSmaller_T_1 : {{1'd0},
    far_alignedSigSmaller}; // @[AddRecFN.scala 97:39]
  wire [13:0] _far_sigSum_T = {far_sigLarger, 3'h0}; // @[AddRecFN.scala 98:36]
  wire [14:0] _GEN_3 = {{1'd0}, _far_sigSum_T}; // @[AddRecFN.scala 98:41]
  wire [14:0] _far_sigSum_T_2 = _GEN_3 + far_negAlignedSigSmaller; // @[AddRecFN.scala 98:41]
  wire [14:0] _GEN_4 = {{14'd0}, _closeSubMags_T}; // @[AddRecFN.scala 98:68]
  wire [14:0] far_sigSum = _far_sigSum_T_2 + _GEN_4; // @[AddRecFN.scala 98:68]
  wire [13:0] _GEN_5 = {{13'd0}, far_sigSum[0]}; // @[AddRecFN.scala 99:67]
  wire [13:0] _far_sigOut_T_2 = far_sigSum[14:1] | _GEN_5; // @[AddRecFN.scala 99:67]
  wire [14:0] _far_sigOut_T_3 = _closeSubMags_T ? far_sigSum : {{1'd0}, _far_sigOut_T_2}; // @[AddRecFN.scala 99:25]
  wire [13:0] far_sigOut = _far_sigOut_T_3[13:0]; // @[AddRecFN.scala 99:83]
  wire  notSigNaN_invalidExc = io_a_isInf & io_b_isInf & _closeSubMags_T; // @[AddRecFN.scala 102:57]
  wire  notNaN_isInfOut = io_a_isInf | io_b_isInf; // @[AddRecFN.scala 103:38]
  wire  addZeros = io_a_isZero & io_b_isZero; // @[AddRecFN.scala 104:32]
  wire  notNaN_specialCase = notNaN_isInfOut | addZeros; // @[AddRecFN.scala 105:46]
  wire  _notNaN_signOut_T_1 = io_a_isInf & io_a_sign; // @[AddRecFN.scala 109:39]
  wire  _notNaN_signOut_T_2 = eqSigns & io_a_sign | _notNaN_signOut_T_1; // @[AddRecFN.scala 108:63]
  wire  _notNaN_signOut_T_3 = io_b_isInf & effSignB; // @[AddRecFN.scala 110:39]
  wire  _notNaN_signOut_T_4 = _notNaN_signOut_T_2 | _notNaN_signOut_T_3; // @[AddRecFN.scala 109:63]
  wire  _notNaN_signOut_T_9 = ~notNaN_specialCase; // @[AddRecFN.scala 112:10]
  wire  _notNaN_signOut_T_12 = ~notNaN_specialCase & closeSubMags & ~close_totalCancellation; // @[AddRecFN.scala 112:46]
  wire  _notNaN_signOut_T_13 = _notNaN_signOut_T_12 & close_notTotalCancellation_signOut; // @[AddRecFN.scala 113:38]
  wire  _notNaN_signOut_T_14 = _notNaN_signOut_T_4 | _notNaN_signOut_T_13; // @[AddRecFN.scala 111:63]
  wire  _notNaN_signOut_T_18 = _notNaN_signOut_T_9 & ~closeSubMags & far_signOut; // @[AddRecFN.scala 114:47]
  wire [6:0] _common_sExpOut_T_2 = closeSubMags | _modNatAlignDist_T ? $signed(io_b_sExp) : $signed(io_a_sExp); // @[AddRecFN.scala 116:13]
  wire [3:0] _common_sExpOut_T_3 = closeSubMags ? close_nearNormDist : {{3'd0}, _closeSubMags_T}; // @[AddRecFN.scala 117:18]
  wire [4:0] _common_sExpOut_T_4 = {1'b0,$signed(_common_sExpOut_T_3)}; // @[AddRecFN.scala 117:66]
  wire [6:0] _GEN_6 = {{2{_common_sExpOut_T_4[4]}},_common_sExpOut_T_4}; // @[AddRecFN.scala 117:13]
  wire  _io_invalidExc_T_2 = io_a_isNaN & ~io_a_sig[9]; // @[common.scala 82:46]
  wire  _io_invalidExc_T_5 = io_b_isNaN & ~io_b_sig[9]; // @[common.scala 82:46]
  assign io_invalidExc = _io_invalidExc_T_2 | _io_invalidExc_T_5 | notSigNaN_invalidExc; // @[AddRecFN.scala 121:71]
  assign io_rawOut_isNaN = io_a_isNaN | io_b_isNaN; // @[AddRecFN.scala 125:35]
  assign io_rawOut_isInf = io_a_isInf | io_b_isInf; // @[AddRecFN.scala 103:38]
  assign io_rawOut_isZero = addZeros | ~notNaN_isInfOut & closeSubMags & close_totalCancellation; // @[AddRecFN.scala 106:37]
  assign io_rawOut_sign = _notNaN_signOut_T_14 | _notNaN_signOut_T_18; // @[AddRecFN.scala 113:77]
  assign io_rawOut_sExp = $signed(_common_sExpOut_T_2) - $signed(_GEN_6); // @[AddRecFN.scala 117:13]
  assign io_rawOut_sig = closeSubMags ? close_sigOut : far_sigOut; // @[AddRecFN.scala 118:28]
endmodule
module RoundAnyRawFNToRecFN(
  input         io_invalidExc,
  input         io_in_isNaN,
  input         io_in_isInf,
  input         io_in_isZero,
  input         io_in_sign,
  input  [6:0]  io_in_sExp,
  input  [13:0] io_in_sig,
  output [16:0] io_out
);
  wire  doShiftSigDown1 = io_in_sig[13]; // @[RoundAnyRawFNToRecFN.scala 118:61]
  wire [5:0] _roundMask_T_1 = ~io_in_sExp[5:0]; // @[primitives.scala 51:21]
  wire [64:0] roundMask_shift = 65'sh10000000000000000 >>> _roundMask_T_1; // @[primitives.scala 77:58]
  wire [7:0] _GEN_0 = {{4'd0}, roundMask_shift[14:11]}; // @[Bitwise.scala 108:31]
  wire [7:0] _roundMask_T_7 = _GEN_0 & 8'hf; // @[Bitwise.scala 108:31]
  wire [7:0] _roundMask_T_9 = {roundMask_shift[10:7], 4'h0}; // @[Bitwise.scala 108:70]
  wire [7:0] _roundMask_T_11 = _roundMask_T_9 & 8'hf0; // @[Bitwise.scala 108:80]
  wire [7:0] _roundMask_T_12 = _roundMask_T_7 | _roundMask_T_11; // @[Bitwise.scala 108:39]
  wire [7:0] _GEN_1 = {{2'd0}, _roundMask_T_12[7:2]}; // @[Bitwise.scala 108:31]
  wire [7:0] _roundMask_T_17 = _GEN_1 & 8'h33; // @[Bitwise.scala 108:31]
  wire [7:0] _roundMask_T_19 = {_roundMask_T_12[5:0], 2'h0}; // @[Bitwise.scala 108:70]
  wire [7:0] _roundMask_T_21 = _roundMask_T_19 & 8'hcc; // @[Bitwise.scala 108:80]
  wire [7:0] _roundMask_T_22 = _roundMask_T_17 | _roundMask_T_21; // @[Bitwise.scala 108:39]
  wire [7:0] _GEN_2 = {{1'd0}, _roundMask_T_22[7:1]}; // @[Bitwise.scala 108:31]
  wire [7:0] _roundMask_T_27 = _GEN_2 & 8'h55; // @[Bitwise.scala 108:31]
  wire [7:0] _roundMask_T_29 = {_roundMask_T_22[6:0], 1'h0}; // @[Bitwise.scala 108:70]
  wire [7:0] _roundMask_T_31 = _roundMask_T_29 & 8'haa; // @[Bitwise.scala 108:80]
  wire [7:0] _roundMask_T_32 = _roundMask_T_27 | _roundMask_T_31; // @[Bitwise.scala 108:39]
  wire [11:0] _roundMask_T_43 = {_roundMask_T_32,roundMask_shift[15],roundMask_shift[16],roundMask_shift[17],
    roundMask_shift[18]}; // @[Cat.scala 33:92]
  wire [11:0] _GEN_3 = {{11'd0}, doShiftSigDown1}; // @[RoundAnyRawFNToRecFN.scala 157:23]
  wire [11:0] _roundMask_T_44 = _roundMask_T_43 | _GEN_3; // @[RoundAnyRawFNToRecFN.scala 157:23]
  wire [13:0] roundMask = {_roundMask_T_44,2'h3}; // @[Cat.scala 33:92]
  wire [13:0] shiftedRoundMask = {1'h0,roundMask[13:1]}; // @[Cat.scala 33:92]
  wire [13:0] _roundPosMask_T = ~shiftedRoundMask; // @[RoundAnyRawFNToRecFN.scala 161:28]
  wire [13:0] roundPosMask = _roundPosMask_T & roundMask; // @[RoundAnyRawFNToRecFN.scala 161:46]
  wire [13:0] _roundPosBit_T = io_in_sig & roundPosMask; // @[RoundAnyRawFNToRecFN.scala 162:40]
  wire  roundPosBit = |_roundPosBit_T; // @[RoundAnyRawFNToRecFN.scala 162:56]
  wire [13:0] _anyRoundExtra_T = io_in_sig & shiftedRoundMask; // @[RoundAnyRawFNToRecFN.scala 163:42]
  wire  anyRoundExtra = |_anyRoundExtra_T; // @[RoundAnyRawFNToRecFN.scala 163:62]
  wire [13:0] _roundedSig_T = io_in_sig | roundMask; // @[RoundAnyRawFNToRecFN.scala 172:32]
  wire [12:0] _roundedSig_T_2 = _roundedSig_T[13:2] + 12'h1; // @[RoundAnyRawFNToRecFN.scala 172:49]
  wire  _roundedSig_T_4 = ~anyRoundExtra; // @[RoundAnyRawFNToRecFN.scala 174:30]
  wire [12:0] _roundedSig_T_7 = roundPosBit & _roundedSig_T_4 ? roundMask[13:1] : 13'h0; // @[RoundAnyRawFNToRecFN.scala 173:25]
  wire [12:0] _roundedSig_T_8 = ~_roundedSig_T_7; // @[RoundAnyRawFNToRecFN.scala 173:21]
  wire [12:0] _roundedSig_T_9 = _roundedSig_T_2 & _roundedSig_T_8; // @[RoundAnyRawFNToRecFN.scala 172:61]
  wire [13:0] _roundedSig_T_10 = ~roundMask; // @[RoundAnyRawFNToRecFN.scala 178:32]
  wire [13:0] _roundedSig_T_11 = io_in_sig & _roundedSig_T_10; // @[RoundAnyRawFNToRecFN.scala 178:30]
  wire [12:0] _roundedSig_T_16 = {{1'd0}, _roundedSig_T_11[13:2]}; // @[RoundAnyRawFNToRecFN.scala 178:47]
  wire [12:0] roundedSig = roundPosBit ? _roundedSig_T_9 : _roundedSig_T_16; // @[RoundAnyRawFNToRecFN.scala 171:16]
  wire [2:0] _sRoundedExp_T_1 = {1'b0,$signed(roundedSig[12:11])}; // @[RoundAnyRawFNToRecFN.scala 183:69]
  wire [6:0] _GEN_4 = {{4{_sRoundedExp_T_1[2]}},_sRoundedExp_T_1}; // @[RoundAnyRawFNToRecFN.scala 183:40]
  wire [7:0] sRoundedExp = $signed(io_in_sExp) + $signed(_GEN_4); // @[RoundAnyRawFNToRecFN.scala 183:40]
  wire [5:0] common_expOut = sRoundedExp[5:0]; // @[RoundAnyRawFNToRecFN.scala 185:37]
  wire [9:0] common_fractOut = doShiftSigDown1 ? roundedSig[10:1] : roundedSig[9:0]; // @[RoundAnyRawFNToRecFN.scala 187:16]
  wire [3:0] _common_overflow_T = sRoundedExp[7:4]; // @[RoundAnyRawFNToRecFN.scala 194:30]
  wire  common_overflow = $signed(_common_overflow_T) >= 4'sh3; // @[RoundAnyRawFNToRecFN.scala 194:50]
  wire  common_totalUnderflow = $signed(sRoundedExp) < 8'sh8; // @[RoundAnyRawFNToRecFN.scala 198:31]
  wire  isNaNOut = io_invalidExc | io_in_isNaN; // @[RoundAnyRawFNToRecFN.scala 233:34]
  wire  commonCase = ~isNaNOut & ~io_in_isInf & ~io_in_isZero; // @[RoundAnyRawFNToRecFN.scala 235:61]
  wire  overflow = commonCase & common_overflow; // @[RoundAnyRawFNToRecFN.scala 236:32]
  wire  notNaN_isInfOut = io_in_isInf | overflow; // @[RoundAnyRawFNToRecFN.scala 246:32]
  wire  signOut = isNaNOut ? 1'h0 : io_in_sign; // @[RoundAnyRawFNToRecFN.scala 248:22]
  wire [5:0] _expOut_T_1 = io_in_isZero | common_totalUnderflow ? 6'h38 : 6'h0; // @[RoundAnyRawFNToRecFN.scala 251:18]
  wire [5:0] _expOut_T_2 = ~_expOut_T_1; // @[RoundAnyRawFNToRecFN.scala 251:14]
  wire [5:0] _expOut_T_3 = common_expOut & _expOut_T_2; // @[RoundAnyRawFNToRecFN.scala 250:24]
  wire [5:0] _expOut_T_11 = notNaN_isInfOut ? 6'h8 : 6'h0; // @[RoundAnyRawFNToRecFN.scala 263:18]
  wire [5:0] _expOut_T_12 = ~_expOut_T_11; // @[RoundAnyRawFNToRecFN.scala 263:14]
  wire [5:0] _expOut_T_13 = _expOut_T_3 & _expOut_T_12; // @[RoundAnyRawFNToRecFN.scala 262:17]
  wire [5:0] _expOut_T_18 = notNaN_isInfOut ? 6'h30 : 6'h0; // @[RoundAnyRawFNToRecFN.scala 275:16]
  wire [5:0] _expOut_T_19 = _expOut_T_13 | _expOut_T_18; // @[RoundAnyRawFNToRecFN.scala 274:15]
  wire [5:0] _expOut_T_20 = isNaNOut ? 6'h38 : 6'h0; // @[RoundAnyRawFNToRecFN.scala 276:16]
  wire [5:0] expOut = _expOut_T_19 | _expOut_T_20; // @[RoundAnyRawFNToRecFN.scala 275:77]
  wire [9:0] _fractOut_T_2 = isNaNOut ? 10'h200 : 10'h0; // @[RoundAnyRawFNToRecFN.scala 279:16]
  wire [9:0] fractOut = isNaNOut | io_in_isZero | common_totalUnderflow ? _fractOut_T_2 : common_fractOut; // @[RoundAnyRawFNToRecFN.scala 278:12]
  wire [6:0] io_out_hi = {signOut,expOut}; // @[Cat.scala 33:92]
  assign io_out = {io_out_hi,fractOut}; // @[Cat.scala 33:92]
endmodule
module RoundRawFNToRecFN(
  input         io_invalidExc,
  input         io_in_isNaN,
  input         io_in_isInf,
  input         io_in_isZero,
  input         io_in_sign,
  input  [6:0]  io_in_sExp,
  input  [13:0] io_in_sig,
  output [16:0] io_out
);
  wire  roundAnyRawFNToRecFN_io_invalidExc; // @[RoundAnyRawFNToRecFN.scala 307:15]
  wire  roundAnyRawFNToRecFN_io_in_isNaN; // @[RoundAnyRawFNToRecFN.scala 307:15]
  wire  roundAnyRawFNToRecFN_io_in_isInf; // @[RoundAnyRawFNToRecFN.scala 307:15]
  wire  roundAnyRawFNToRecFN_io_in_isZero; // @[RoundAnyRawFNToRecFN.scala 307:15]
  wire  roundAnyRawFNToRecFN_io_in_sign; // @[RoundAnyRawFNToRecFN.scala 307:15]
  wire [6:0] roundAnyRawFNToRecFN_io_in_sExp; // @[RoundAnyRawFNToRecFN.scala 307:15]
  wire [13:0] roundAnyRawFNToRecFN_io_in_sig; // @[RoundAnyRawFNToRecFN.scala 307:15]
  wire [16:0] roundAnyRawFNToRecFN_io_out; // @[RoundAnyRawFNToRecFN.scala 307:15]
  RoundAnyRawFNToRecFN roundAnyRawFNToRecFN ( // @[RoundAnyRawFNToRecFN.scala 307:15]
    .io_invalidExc(roundAnyRawFNToRecFN_io_invalidExc),
    .io_in_isNaN(roundAnyRawFNToRecFN_io_in_isNaN),
    .io_in_isInf(roundAnyRawFNToRecFN_io_in_isInf),
    .io_in_isZero(roundAnyRawFNToRecFN_io_in_isZero),
    .io_in_sign(roundAnyRawFNToRecFN_io_in_sign),
    .io_in_sExp(roundAnyRawFNToRecFN_io_in_sExp),
    .io_in_sig(roundAnyRawFNToRecFN_io_in_sig),
    .io_out(roundAnyRawFNToRecFN_io_out)
  );
  assign io_out = roundAnyRawFNToRecFN_io_out; // @[RoundAnyRawFNToRecFN.scala 315:23]
  assign roundAnyRawFNToRecFN_io_invalidExc = io_invalidExc; // @[RoundAnyRawFNToRecFN.scala 310:44]
  assign roundAnyRawFNToRecFN_io_in_isNaN = io_in_isNaN; // @[RoundAnyRawFNToRecFN.scala 312:44]
  assign roundAnyRawFNToRecFN_io_in_isInf = io_in_isInf; // @[RoundAnyRawFNToRecFN.scala 312:44]
  assign roundAnyRawFNToRecFN_io_in_isZero = io_in_isZero; // @[RoundAnyRawFNToRecFN.scala 312:44]
  assign roundAnyRawFNToRecFN_io_in_sign = io_in_sign; // @[RoundAnyRawFNToRecFN.scala 312:44]
  assign roundAnyRawFNToRecFN_io_in_sExp = io_in_sExp; // @[RoundAnyRawFNToRecFN.scala 312:44]
  assign roundAnyRawFNToRecFN_io_in_sig = io_in_sig; // @[RoundAnyRawFNToRecFN.scala 312:44]
endmodule
module AddRecFN(
  input         io_subOp,
  input  [16:0] io_a,
  input  [16:0] io_b,
  output [16:0] io_out
);
  wire  addRawFN__io_subOp; // @[AddRecFN.scala 147:26]
  wire  addRawFN__io_a_isNaN; // @[AddRecFN.scala 147:26]
  wire  addRawFN__io_a_isInf; // @[AddRecFN.scala 147:26]
  wire  addRawFN__io_a_isZero; // @[AddRecFN.scala 147:26]
  wire  addRawFN__io_a_sign; // @[AddRecFN.scala 147:26]
  wire [6:0] addRawFN__io_a_sExp; // @[AddRecFN.scala 147:26]
  wire [11:0] addRawFN__io_a_sig; // @[AddRecFN.scala 147:26]
  wire  addRawFN__io_b_isNaN; // @[AddRecFN.scala 147:26]
  wire  addRawFN__io_b_isInf; // @[AddRecFN.scala 147:26]
  wire  addRawFN__io_b_isZero; // @[AddRecFN.scala 147:26]
  wire  addRawFN__io_b_sign; // @[AddRecFN.scala 147:26]
  wire [6:0] addRawFN__io_b_sExp; // @[AddRecFN.scala 147:26]
  wire [11:0] addRawFN__io_b_sig; // @[AddRecFN.scala 147:26]
  wire  addRawFN__io_invalidExc; // @[AddRecFN.scala 147:26]
  wire  addRawFN__io_rawOut_isNaN; // @[AddRecFN.scala 147:26]
  wire  addRawFN__io_rawOut_isInf; // @[AddRecFN.scala 147:26]
  wire  addRawFN__io_rawOut_isZero; // @[AddRecFN.scala 147:26]
  wire  addRawFN__io_rawOut_sign; // @[AddRecFN.scala 147:26]
  wire [6:0] addRawFN__io_rawOut_sExp; // @[AddRecFN.scala 147:26]
  wire [13:0] addRawFN__io_rawOut_sig; // @[AddRecFN.scala 147:26]
  wire  roundRawFNToRecFN_io_invalidExc; // @[AddRecFN.scala 157:15]
  wire  roundRawFNToRecFN_io_in_isNaN; // @[AddRecFN.scala 157:15]
  wire  roundRawFNToRecFN_io_in_isInf; // @[AddRecFN.scala 157:15]
  wire  roundRawFNToRecFN_io_in_isZero; // @[AddRecFN.scala 157:15]
  wire  roundRawFNToRecFN_io_in_sign; // @[AddRecFN.scala 157:15]
  wire [6:0] roundRawFNToRecFN_io_in_sExp; // @[AddRecFN.scala 157:15]
  wire [13:0] roundRawFNToRecFN_io_in_sig; // @[AddRecFN.scala 157:15]
  wire [16:0] roundRawFNToRecFN_io_out; // @[AddRecFN.scala 157:15]
  wire [5:0] addRawFN_io_a_exp = io_a[15:10]; // @[rawFloatFromRecFN.scala 50:21]
  wire  addRawFN_io_a_isZero = addRawFN_io_a_exp[5:3] == 3'h0; // @[rawFloatFromRecFN.scala 51:54]
  wire  addRawFN_io_a_isSpecial = addRawFN_io_a_exp[5:4] == 2'h3; // @[rawFloatFromRecFN.scala 52:54]
  wire  _addRawFN_io_a_out_sig_T = ~addRawFN_io_a_isZero; // @[rawFloatFromRecFN.scala 60:39]
  wire [1:0] addRawFN_io_a_out_sig_hi = {1'h0,_addRawFN_io_a_out_sig_T}; // @[Cat.scala 33:92]
  wire [5:0] addRawFN_io_b_exp = io_b[15:10]; // @[rawFloatFromRecFN.scala 50:21]
  wire  addRawFN_io_b_isZero = addRawFN_io_b_exp[5:3] == 3'h0; // @[rawFloatFromRecFN.scala 51:54]
  wire  addRawFN_io_b_isSpecial = addRawFN_io_b_exp[5:4] == 2'h3; // @[rawFloatFromRecFN.scala 52:54]
  wire  _addRawFN_io_b_out_sig_T = ~addRawFN_io_b_isZero; // @[rawFloatFromRecFN.scala 60:39]
  wire [1:0] addRawFN_io_b_out_sig_hi = {1'h0,_addRawFN_io_b_out_sig_T}; // @[Cat.scala 33:92]
  AddRawFN addRawFN_ ( // @[AddRecFN.scala 147:26]
    .io_subOp(addRawFN__io_subOp),
    .io_a_isNaN(addRawFN__io_a_isNaN),
    .io_a_isInf(addRawFN__io_a_isInf),
    .io_a_isZero(addRawFN__io_a_isZero),
    .io_a_sign(addRawFN__io_a_sign),
    .io_a_sExp(addRawFN__io_a_sExp),
    .io_a_sig(addRawFN__io_a_sig),
    .io_b_isNaN(addRawFN__io_b_isNaN),
    .io_b_isInf(addRawFN__io_b_isInf),
    .io_b_isZero(addRawFN__io_b_isZero),
    .io_b_sign(addRawFN__io_b_sign),
    .io_b_sExp(addRawFN__io_b_sExp),
    .io_b_sig(addRawFN__io_b_sig),
    .io_invalidExc(addRawFN__io_invalidExc),
    .io_rawOut_isNaN(addRawFN__io_rawOut_isNaN),
    .io_rawOut_isInf(addRawFN__io_rawOut_isInf),
    .io_rawOut_isZero(addRawFN__io_rawOut_isZero),
    .io_rawOut_sign(addRawFN__io_rawOut_sign),
    .io_rawOut_sExp(addRawFN__io_rawOut_sExp),
    .io_rawOut_sig(addRawFN__io_rawOut_sig)
  );
  RoundRawFNToRecFN roundRawFNToRecFN ( // @[AddRecFN.scala 157:15]
    .io_invalidExc(roundRawFNToRecFN_io_invalidExc),
    .io_in_isNaN(roundRawFNToRecFN_io_in_isNaN),
    .io_in_isInf(roundRawFNToRecFN_io_in_isInf),
    .io_in_isZero(roundRawFNToRecFN_io_in_isZero),
    .io_in_sign(roundRawFNToRecFN_io_in_sign),
    .io_in_sExp(roundRawFNToRecFN_io_in_sExp),
    .io_in_sig(roundRawFNToRecFN_io_in_sig),
    .io_out(roundRawFNToRecFN_io_out)
  );
  assign io_out = roundRawFNToRecFN_io_out; // @[AddRecFN.scala 163:23]
  assign addRawFN__io_subOp = io_subOp; // @[AddRecFN.scala 149:30]
  assign addRawFN__io_a_isNaN = addRawFN_io_a_isSpecial & addRawFN_io_a_exp[3]; // @[rawFloatFromRecFN.scala 55:33]
  assign addRawFN__io_a_isInf = addRawFN_io_a_isSpecial & ~addRawFN_io_a_exp[3]; // @[rawFloatFromRecFN.scala 56:33]
  assign addRawFN__io_a_isZero = addRawFN_io_a_exp[5:3] == 3'h0; // @[rawFloatFromRecFN.scala 51:54]
  assign addRawFN__io_a_sign = io_a[16]; // @[rawFloatFromRecFN.scala 58:25]
  assign addRawFN__io_a_sExp = {1'b0,$signed(addRawFN_io_a_exp)}; // @[rawFloatFromRecFN.scala 59:27]
  assign addRawFN__io_a_sig = {addRawFN_io_a_out_sig_hi,io_a[9:0]}; // @[Cat.scala 33:92]
  assign addRawFN__io_b_isNaN = addRawFN_io_b_isSpecial & addRawFN_io_b_exp[3]; // @[rawFloatFromRecFN.scala 55:33]
  assign addRawFN__io_b_isInf = addRawFN_io_b_isSpecial & ~addRawFN_io_b_exp[3]; // @[rawFloatFromRecFN.scala 56:33]
  assign addRawFN__io_b_isZero = addRawFN_io_b_exp[5:3] == 3'h0; // @[rawFloatFromRecFN.scala 51:54]
  assign addRawFN__io_b_sign = io_b[16]; // @[rawFloatFromRecFN.scala 58:25]
  assign addRawFN__io_b_sExp = {1'b0,$signed(addRawFN_io_b_exp)}; // @[rawFloatFromRecFN.scala 59:27]
  assign addRawFN__io_b_sig = {addRawFN_io_b_out_sig_hi,io_b[9:0]}; // @[Cat.scala 33:92]
  assign roundRawFNToRecFN_io_invalidExc = addRawFN__io_invalidExc; // @[AddRecFN.scala 158:39]
  assign roundRawFNToRecFN_io_in_isNaN = addRawFN__io_rawOut_isNaN; // @[AddRecFN.scala 160:39]
  assign roundRawFNToRecFN_io_in_isInf = addRawFN__io_rawOut_isInf; // @[AddRecFN.scala 160:39]
  assign roundRawFNToRecFN_io_in_isZero = addRawFN__io_rawOut_isZero; // @[AddRecFN.scala 160:39]
  assign roundRawFNToRecFN_io_in_sign = addRawFN__io_rawOut_sign; // @[AddRecFN.scala 160:39]
  assign roundRawFNToRecFN_io_in_sExp = addRawFN__io_rawOut_sExp; // @[AddRecFN.scala 160:39]
  assign roundRawFNToRecFN_io_in_sig = addRawFN__io_rawOut_sig; // @[AddRecFN.scala 160:39]
endmodule
module FloatAdd(
  input  [16:0] io_op1,
  input  [16:0] io_op2,
  output [16:0] io_res
);
  wire  float_adder_io_subOp; // @[Float.scala 14:27]
  wire [16:0] float_adder_io_a; // @[Float.scala 14:27]
  wire [16:0] float_adder_io_b; // @[Float.scala 14:27]
  wire [16:0] float_adder_io_out; // @[Float.scala 14:27]
  AddRecFN float_adder ( // @[Float.scala 14:27]
    .io_subOp(float_adder_io_subOp),
    .io_a(float_adder_io_a),
    .io_b(float_adder_io_b),
    .io_out(float_adder_io_out)
  );
  assign io_res = float_adder_io_out; // @[Float.scala 20:10]
  assign float_adder_io_subOp = 1'h0; // @[Float.scala 15:24]
  assign float_adder_io_a = io_op1; // @[Float.scala 16:20]
  assign float_adder_io_b = io_op2; // @[Float.scala 17:20]
endmodule
module ComplexAdd(
  input  [16:0] io_op1_re,
  input  [16:0] io_op1_im,
  input  [16:0] io_op2_re,
  input  [16:0] io_op2_im,
  output [16:0] io_res_re,
  output [16:0] io_res_im
);
  wire [16:0] io_res_re_inst_io_op1; // @[Float.scala 25:22]
  wire [16:0] io_res_re_inst_io_op2; // @[Float.scala 25:22]
  wire [16:0] io_res_re_inst_io_res; // @[Float.scala 25:22]
  wire [16:0] io_res_im_inst_io_op1; // @[Float.scala 25:22]
  wire [16:0] io_res_im_inst_io_op2; // @[Float.scala 25:22]
  wire [16:0] io_res_im_inst_io_res; // @[Float.scala 25:22]
  FloatAdd io_res_re_inst ( // @[Float.scala 25:22]
    .io_op1(io_res_re_inst_io_op1),
    .io_op2(io_res_re_inst_io_op2),
    .io_res(io_res_re_inst_io_res)
  );
  FloatAdd io_res_im_inst ( // @[Float.scala 25:22]
    .io_op1(io_res_im_inst_io_op1),
    .io_op2(io_res_im_inst_io_op2),
    .io_res(io_res_im_inst_io_res)
  );
  assign io_res_re = io_res_re_inst_io_res; // @[Modules.scala 71:15]
  assign io_res_im = io_res_im_inst_io_res; // @[Modules.scala 72:15]
  assign io_res_re_inst_io_op1 = io_op1_re; // @[Float.scala 26:17]
  assign io_res_re_inst_io_op2 = io_op2_re; // @[Float.scala 27:17]
  assign io_res_im_inst_io_op1 = io_op1_im; // @[Float.scala 26:17]
  assign io_res_im_inst_io_op2 = io_op2_im; // @[Float.scala 27:17]
endmodule
module FloatSub(
  input  [16:0] io_op1,
  input  [16:0] io_op2,
  output [16:0] io_res
);
  wire  float_adder_io_subOp; // @[Float.scala 34:27]
  wire [16:0] float_adder_io_a; // @[Float.scala 34:27]
  wire [16:0] float_adder_io_b; // @[Float.scala 34:27]
  wire [16:0] float_adder_io_out; // @[Float.scala 34:27]
  AddRecFN float_adder ( // @[Float.scala 34:27]
    .io_subOp(float_adder_io_subOp),
    .io_a(float_adder_io_a),
    .io_b(float_adder_io_b),
    .io_out(float_adder_io_out)
  );
  assign io_res = float_adder_io_out; // @[Float.scala 40:10]
  assign float_adder_io_subOp = 1'h1; // @[Float.scala 35:24]
  assign float_adder_io_a = io_op1; // @[Float.scala 36:20]
  assign float_adder_io_b = io_op2; // @[Float.scala 37:20]
endmodule
module ComplexSub(
  input  [16:0] io_op1_re,
  input  [16:0] io_op1_im,
  input  [16:0] io_op2_re,
  input  [16:0] io_op2_im,
  output [16:0] io_res_re,
  output [16:0] io_res_im
);
  wire [16:0] io_res_re_inst_io_op1; // @[Float.scala 45:22]
  wire [16:0] io_res_re_inst_io_op2; // @[Float.scala 45:22]
  wire [16:0] io_res_re_inst_io_res; // @[Float.scala 45:22]
  wire [16:0] io_res_im_inst_io_op1; // @[Float.scala 45:22]
  wire [16:0] io_res_im_inst_io_op2; // @[Float.scala 45:22]
  wire [16:0] io_res_im_inst_io_res; // @[Float.scala 45:22]
  FloatSub io_res_re_inst ( // @[Float.scala 45:22]
    .io_op1(io_res_re_inst_io_op1),
    .io_op2(io_res_re_inst_io_op2),
    .io_res(io_res_re_inst_io_res)
  );
  FloatSub io_res_im_inst ( // @[Float.scala 45:22]
    .io_op1(io_res_im_inst_io_op1),
    .io_op2(io_res_im_inst_io_op2),
    .io_res(io_res_im_inst_io_res)
  );
  assign io_res_re = io_res_re_inst_io_res; // @[Modules.scala 90:15]
  assign io_res_im = io_res_im_inst_io_res; // @[Modules.scala 91:15]
  assign io_res_re_inst_io_op1 = io_op1_re; // @[Float.scala 46:17]
  assign io_res_re_inst_io_op2 = io_op2_re; // @[Float.scala 47:17]
  assign io_res_im_inst_io_op1 = io_op1_im; // @[Float.scala 46:17]
  assign io_res_im_inst_io_op2 = io_op2_im; // @[Float.scala 47:17]
endmodule
module MulFullRawFN(
  input         io_a_isNaN,
  input         io_a_isInf,
  input         io_a_isZero,
  input         io_a_sign,
  input  [6:0]  io_a_sExp,
  input  [11:0] io_a_sig,
  input         io_b_isNaN,
  input         io_b_isInf,
  input         io_b_isZero,
  input         io_b_sign,
  input  [6:0]  io_b_sExp,
  input  [11:0] io_b_sig,
  output        io_invalidExc,
  output        io_rawOut_isNaN,
  output        io_rawOut_isInf,
  output        io_rawOut_isZero,
  output        io_rawOut_sign,
  output [6:0]  io_rawOut_sExp,
  output [21:0] io_rawOut_sig
);
  wire  notSigNaN_invalidExc = io_a_isInf & io_b_isZero | io_a_isZero & io_b_isInf; // @[MulRecFN.scala 58:60]
  wire [6:0] _common_sExpOut_T_2 = $signed(io_a_sExp) + $signed(io_b_sExp); // @[MulRecFN.scala 62:36]
  wire [23:0] _common_sigOut_T = io_a_sig * io_b_sig; // @[MulRecFN.scala 63:35]
  wire  _io_invalidExc_T_2 = io_a_isNaN & ~io_a_sig[9]; // @[common.scala 82:46]
  wire  _io_invalidExc_T_5 = io_b_isNaN & ~io_b_sig[9]; // @[common.scala 82:46]
  assign io_invalidExc = _io_invalidExc_T_2 | _io_invalidExc_T_5 | notSigNaN_invalidExc; // @[MulRecFN.scala 66:71]
  assign io_rawOut_isNaN = io_a_isNaN | io_b_isNaN; // @[MulRecFN.scala 70:35]
  assign io_rawOut_isInf = io_a_isInf | io_b_isInf; // @[MulRecFN.scala 59:38]
  assign io_rawOut_isZero = io_a_isZero | io_b_isZero; // @[MulRecFN.scala 60:40]
  assign io_rawOut_sign = io_a_sign ^ io_b_sign; // @[MulRecFN.scala 61:36]
  assign io_rawOut_sExp = $signed(_common_sExpOut_T_2) - 7'sh20; // @[MulRecFN.scala 62:48]
  assign io_rawOut_sig = _common_sigOut_T[21:0]; // @[MulRecFN.scala 63:46]
endmodule
module MulRawFN(
  input         io_a_isNaN,
  input         io_a_isInf,
  input         io_a_isZero,
  input         io_a_sign,
  input  [6:0]  io_a_sExp,
  input  [11:0] io_a_sig,
  input         io_b_isNaN,
  input         io_b_isInf,
  input         io_b_isZero,
  input         io_b_sign,
  input  [6:0]  io_b_sExp,
  input  [11:0] io_b_sig,
  output        io_invalidExc,
  output        io_rawOut_isNaN,
  output        io_rawOut_isInf,
  output        io_rawOut_isZero,
  output        io_rawOut_sign,
  output [6:0]  io_rawOut_sExp,
  output [13:0] io_rawOut_sig
);
  wire  mulFullRaw_io_a_isNaN; // @[MulRecFN.scala 84:28]
  wire  mulFullRaw_io_a_isInf; // @[MulRecFN.scala 84:28]
  wire  mulFullRaw_io_a_isZero; // @[MulRecFN.scala 84:28]
  wire  mulFullRaw_io_a_sign; // @[MulRecFN.scala 84:28]
  wire [6:0] mulFullRaw_io_a_sExp; // @[MulRecFN.scala 84:28]
  wire [11:0] mulFullRaw_io_a_sig; // @[MulRecFN.scala 84:28]
  wire  mulFullRaw_io_b_isNaN; // @[MulRecFN.scala 84:28]
  wire  mulFullRaw_io_b_isInf; // @[MulRecFN.scala 84:28]
  wire  mulFullRaw_io_b_isZero; // @[MulRecFN.scala 84:28]
  wire  mulFullRaw_io_b_sign; // @[MulRecFN.scala 84:28]
  wire [6:0] mulFullRaw_io_b_sExp; // @[MulRecFN.scala 84:28]
  wire [11:0] mulFullRaw_io_b_sig; // @[MulRecFN.scala 84:28]
  wire  mulFullRaw_io_invalidExc; // @[MulRecFN.scala 84:28]
  wire  mulFullRaw_io_rawOut_isNaN; // @[MulRecFN.scala 84:28]
  wire  mulFullRaw_io_rawOut_isInf; // @[MulRecFN.scala 84:28]
  wire  mulFullRaw_io_rawOut_isZero; // @[MulRecFN.scala 84:28]
  wire  mulFullRaw_io_rawOut_sign; // @[MulRecFN.scala 84:28]
  wire [6:0] mulFullRaw_io_rawOut_sExp; // @[MulRecFN.scala 84:28]
  wire [21:0] mulFullRaw_io_rawOut_sig; // @[MulRecFN.scala 84:28]
  wire  _io_rawOut_sig_T_2 = |mulFullRaw_io_rawOut_sig[8:0]; // @[MulRecFN.scala 93:55]
  MulFullRawFN mulFullRaw ( // @[MulRecFN.scala 84:28]
    .io_a_isNaN(mulFullRaw_io_a_isNaN),
    .io_a_isInf(mulFullRaw_io_a_isInf),
    .io_a_isZero(mulFullRaw_io_a_isZero),
    .io_a_sign(mulFullRaw_io_a_sign),
    .io_a_sExp(mulFullRaw_io_a_sExp),
    .io_a_sig(mulFullRaw_io_a_sig),
    .io_b_isNaN(mulFullRaw_io_b_isNaN),
    .io_b_isInf(mulFullRaw_io_b_isInf),
    .io_b_isZero(mulFullRaw_io_b_isZero),
    .io_b_sign(mulFullRaw_io_b_sign),
    .io_b_sExp(mulFullRaw_io_b_sExp),
    .io_b_sig(mulFullRaw_io_b_sig),
    .io_invalidExc(mulFullRaw_io_invalidExc),
    .io_rawOut_isNaN(mulFullRaw_io_rawOut_isNaN),
    .io_rawOut_isInf(mulFullRaw_io_rawOut_isInf),
    .io_rawOut_isZero(mulFullRaw_io_rawOut_isZero),
    .io_rawOut_sign(mulFullRaw_io_rawOut_sign),
    .io_rawOut_sExp(mulFullRaw_io_rawOut_sExp),
    .io_rawOut_sig(mulFullRaw_io_rawOut_sig)
  );
  assign io_invalidExc = mulFullRaw_io_invalidExc; // @[MulRecFN.scala 89:19]
  assign io_rawOut_isNaN = mulFullRaw_io_rawOut_isNaN; // @[MulRecFN.scala 90:15]
  assign io_rawOut_isInf = mulFullRaw_io_rawOut_isInf; // @[MulRecFN.scala 90:15]
  assign io_rawOut_isZero = mulFullRaw_io_rawOut_isZero; // @[MulRecFN.scala 90:15]
  assign io_rawOut_sign = mulFullRaw_io_rawOut_sign; // @[MulRecFN.scala 90:15]
  assign io_rawOut_sExp = mulFullRaw_io_rawOut_sExp; // @[MulRecFN.scala 90:15]
  assign io_rawOut_sig = {mulFullRaw_io_rawOut_sig[21:9],_io_rawOut_sig_T_2}; // @[Cat.scala 33:92]
  assign mulFullRaw_io_a_isNaN = io_a_isNaN; // @[MulRecFN.scala 86:21]
  assign mulFullRaw_io_a_isInf = io_a_isInf; // @[MulRecFN.scala 86:21]
  assign mulFullRaw_io_a_isZero = io_a_isZero; // @[MulRecFN.scala 86:21]
  assign mulFullRaw_io_a_sign = io_a_sign; // @[MulRecFN.scala 86:21]
  assign mulFullRaw_io_a_sExp = io_a_sExp; // @[MulRecFN.scala 86:21]
  assign mulFullRaw_io_a_sig = io_a_sig; // @[MulRecFN.scala 86:21]
  assign mulFullRaw_io_b_isNaN = io_b_isNaN; // @[MulRecFN.scala 87:21]
  assign mulFullRaw_io_b_isInf = io_b_isInf; // @[MulRecFN.scala 87:21]
  assign mulFullRaw_io_b_isZero = io_b_isZero; // @[MulRecFN.scala 87:21]
  assign mulFullRaw_io_b_sign = io_b_sign; // @[MulRecFN.scala 87:21]
  assign mulFullRaw_io_b_sExp = io_b_sExp; // @[MulRecFN.scala 87:21]
  assign mulFullRaw_io_b_sig = io_b_sig; // @[MulRecFN.scala 87:21]
endmodule
module MulRecFN(
  input  [16:0] io_a,
  input  [16:0] io_b,
  output [16:0] io_out
);
  wire  mulRawFN__io_a_isNaN; // @[MulRecFN.scala 113:26]
  wire  mulRawFN__io_a_isInf; // @[MulRecFN.scala 113:26]
  wire  mulRawFN__io_a_isZero; // @[MulRecFN.scala 113:26]
  wire  mulRawFN__io_a_sign; // @[MulRecFN.scala 113:26]
  wire [6:0] mulRawFN__io_a_sExp; // @[MulRecFN.scala 113:26]
  wire [11:0] mulRawFN__io_a_sig; // @[MulRecFN.scala 113:26]
  wire  mulRawFN__io_b_isNaN; // @[MulRecFN.scala 113:26]
  wire  mulRawFN__io_b_isInf; // @[MulRecFN.scala 113:26]
  wire  mulRawFN__io_b_isZero; // @[MulRecFN.scala 113:26]
  wire  mulRawFN__io_b_sign; // @[MulRecFN.scala 113:26]
  wire [6:0] mulRawFN__io_b_sExp; // @[MulRecFN.scala 113:26]
  wire [11:0] mulRawFN__io_b_sig; // @[MulRecFN.scala 113:26]
  wire  mulRawFN__io_invalidExc; // @[MulRecFN.scala 113:26]
  wire  mulRawFN__io_rawOut_isNaN; // @[MulRecFN.scala 113:26]
  wire  mulRawFN__io_rawOut_isInf; // @[MulRecFN.scala 113:26]
  wire  mulRawFN__io_rawOut_isZero; // @[MulRecFN.scala 113:26]
  wire  mulRawFN__io_rawOut_sign; // @[MulRecFN.scala 113:26]
  wire [6:0] mulRawFN__io_rawOut_sExp; // @[MulRecFN.scala 113:26]
  wire [13:0] mulRawFN__io_rawOut_sig; // @[MulRecFN.scala 113:26]
  wire  roundRawFNToRecFN_io_invalidExc; // @[MulRecFN.scala 121:15]
  wire  roundRawFNToRecFN_io_in_isNaN; // @[MulRecFN.scala 121:15]
  wire  roundRawFNToRecFN_io_in_isInf; // @[MulRecFN.scala 121:15]
  wire  roundRawFNToRecFN_io_in_isZero; // @[MulRecFN.scala 121:15]
  wire  roundRawFNToRecFN_io_in_sign; // @[MulRecFN.scala 121:15]
  wire [6:0] roundRawFNToRecFN_io_in_sExp; // @[MulRecFN.scala 121:15]
  wire [13:0] roundRawFNToRecFN_io_in_sig; // @[MulRecFN.scala 121:15]
  wire [16:0] roundRawFNToRecFN_io_out; // @[MulRecFN.scala 121:15]
  wire [5:0] mulRawFN_io_a_exp = io_a[15:10]; // @[rawFloatFromRecFN.scala 50:21]
  wire  mulRawFN_io_a_isZero = mulRawFN_io_a_exp[5:3] == 3'h0; // @[rawFloatFromRecFN.scala 51:54]
  wire  mulRawFN_io_a_isSpecial = mulRawFN_io_a_exp[5:4] == 2'h3; // @[rawFloatFromRecFN.scala 52:54]
  wire  _mulRawFN_io_a_out_sig_T = ~mulRawFN_io_a_isZero; // @[rawFloatFromRecFN.scala 60:39]
  wire [1:0] mulRawFN_io_a_out_sig_hi = {1'h0,_mulRawFN_io_a_out_sig_T}; // @[Cat.scala 33:92]
  wire [5:0] mulRawFN_io_b_exp = io_b[15:10]; // @[rawFloatFromRecFN.scala 50:21]
  wire  mulRawFN_io_b_isZero = mulRawFN_io_b_exp[5:3] == 3'h0; // @[rawFloatFromRecFN.scala 51:54]
  wire  mulRawFN_io_b_isSpecial = mulRawFN_io_b_exp[5:4] == 2'h3; // @[rawFloatFromRecFN.scala 52:54]
  wire  _mulRawFN_io_b_out_sig_T = ~mulRawFN_io_b_isZero; // @[rawFloatFromRecFN.scala 60:39]
  wire [1:0] mulRawFN_io_b_out_sig_hi = {1'h0,_mulRawFN_io_b_out_sig_T}; // @[Cat.scala 33:92]
  MulRawFN mulRawFN_ ( // @[MulRecFN.scala 113:26]
    .io_a_isNaN(mulRawFN__io_a_isNaN),
    .io_a_isInf(mulRawFN__io_a_isInf),
    .io_a_isZero(mulRawFN__io_a_isZero),
    .io_a_sign(mulRawFN__io_a_sign),
    .io_a_sExp(mulRawFN__io_a_sExp),
    .io_a_sig(mulRawFN__io_a_sig),
    .io_b_isNaN(mulRawFN__io_b_isNaN),
    .io_b_isInf(mulRawFN__io_b_isInf),
    .io_b_isZero(mulRawFN__io_b_isZero),
    .io_b_sign(mulRawFN__io_b_sign),
    .io_b_sExp(mulRawFN__io_b_sExp),
    .io_b_sig(mulRawFN__io_b_sig),
    .io_invalidExc(mulRawFN__io_invalidExc),
    .io_rawOut_isNaN(mulRawFN__io_rawOut_isNaN),
    .io_rawOut_isInf(mulRawFN__io_rawOut_isInf),
    .io_rawOut_isZero(mulRawFN__io_rawOut_isZero),
    .io_rawOut_sign(mulRawFN__io_rawOut_sign),
    .io_rawOut_sExp(mulRawFN__io_rawOut_sExp),
    .io_rawOut_sig(mulRawFN__io_rawOut_sig)
  );
  RoundRawFNToRecFN roundRawFNToRecFN ( // @[MulRecFN.scala 121:15]
    .io_invalidExc(roundRawFNToRecFN_io_invalidExc),
    .io_in_isNaN(roundRawFNToRecFN_io_in_isNaN),
    .io_in_isInf(roundRawFNToRecFN_io_in_isInf),
    .io_in_isZero(roundRawFNToRecFN_io_in_isZero),
    .io_in_sign(roundRawFNToRecFN_io_in_sign),
    .io_in_sExp(roundRawFNToRecFN_io_in_sExp),
    .io_in_sig(roundRawFNToRecFN_io_in_sig),
    .io_out(roundRawFNToRecFN_io_out)
  );
  assign io_out = roundRawFNToRecFN_io_out; // @[MulRecFN.scala 127:23]
  assign mulRawFN__io_a_isNaN = mulRawFN_io_a_isSpecial & mulRawFN_io_a_exp[3]; // @[rawFloatFromRecFN.scala 55:33]
  assign mulRawFN__io_a_isInf = mulRawFN_io_a_isSpecial & ~mulRawFN_io_a_exp[3]; // @[rawFloatFromRecFN.scala 56:33]
  assign mulRawFN__io_a_isZero = mulRawFN_io_a_exp[5:3] == 3'h0; // @[rawFloatFromRecFN.scala 51:54]
  assign mulRawFN__io_a_sign = io_a[16]; // @[rawFloatFromRecFN.scala 58:25]
  assign mulRawFN__io_a_sExp = {1'b0,$signed(mulRawFN_io_a_exp)}; // @[rawFloatFromRecFN.scala 59:27]
  assign mulRawFN__io_a_sig = {mulRawFN_io_a_out_sig_hi,io_a[9:0]}; // @[Cat.scala 33:92]
  assign mulRawFN__io_b_isNaN = mulRawFN_io_b_isSpecial & mulRawFN_io_b_exp[3]; // @[rawFloatFromRecFN.scala 55:33]
  assign mulRawFN__io_b_isInf = mulRawFN_io_b_isSpecial & ~mulRawFN_io_b_exp[3]; // @[rawFloatFromRecFN.scala 56:33]
  assign mulRawFN__io_b_isZero = mulRawFN_io_b_exp[5:3] == 3'h0; // @[rawFloatFromRecFN.scala 51:54]
  assign mulRawFN__io_b_sign = io_b[16]; // @[rawFloatFromRecFN.scala 58:25]
  assign mulRawFN__io_b_sExp = {1'b0,$signed(mulRawFN_io_b_exp)}; // @[rawFloatFromRecFN.scala 59:27]
  assign mulRawFN__io_b_sig = {mulRawFN_io_b_out_sig_hi,io_b[9:0]}; // @[Cat.scala 33:92]
  assign roundRawFNToRecFN_io_invalidExc = mulRawFN__io_invalidExc; // @[MulRecFN.scala 122:39]
  assign roundRawFNToRecFN_io_in_isNaN = mulRawFN__io_rawOut_isNaN; // @[MulRecFN.scala 124:39]
  assign roundRawFNToRecFN_io_in_isInf = mulRawFN__io_rawOut_isInf; // @[MulRecFN.scala 124:39]
  assign roundRawFNToRecFN_io_in_isZero = mulRawFN__io_rawOut_isZero; // @[MulRecFN.scala 124:39]
  assign roundRawFNToRecFN_io_in_sign = mulRawFN__io_rawOut_sign; // @[MulRecFN.scala 124:39]
  assign roundRawFNToRecFN_io_in_sExp = mulRawFN__io_rawOut_sExp; // @[MulRecFN.scala 124:39]
  assign roundRawFNToRecFN_io_in_sig = mulRawFN__io_rawOut_sig; // @[MulRecFN.scala 124:39]
endmodule
module FloatMul(
  input  [16:0] io_op1,
  input  [16:0] io_op2,
  output [16:0] io_res
);
  wire [16:0] float_adder_io_a; // @[Float.scala 54:27]
  wire [16:0] float_adder_io_b; // @[Float.scala 54:27]
  wire [16:0] float_adder_io_out; // @[Float.scala 54:27]
  MulRecFN float_adder ( // @[Float.scala 54:27]
    .io_a(float_adder_io_a),
    .io_b(float_adder_io_b),
    .io_out(float_adder_io_out)
  );
  assign io_res = float_adder_io_out; // @[Float.scala 59:10]
  assign float_adder_io_a = io_op1; // @[Float.scala 55:20]
  assign float_adder_io_b = io_op2; // @[Float.scala 56:20]
endmodule
module ComplexMul(
  input  [16:0] io_op1_re,
  input  [16:0] io_op1_im,
  input  [16:0] io_op2_re,
  input  [16:0] io_op2_im,
  output [16:0] io_res_re,
  output [16:0] io_res_im
);
  wire [16:0] io_res_re_inst_io_op1; // @[Float.scala 64:22]
  wire [16:0] io_res_re_inst_io_op2; // @[Float.scala 64:22]
  wire [16:0] io_res_re_inst_io_res; // @[Float.scala 64:22]
  wire [16:0] io_res_re_inst_1_io_op1; // @[Float.scala 64:22]
  wire [16:0] io_res_re_inst_1_io_op2; // @[Float.scala 64:22]
  wire [16:0] io_res_re_inst_1_io_res; // @[Float.scala 64:22]
  wire [16:0] io_res_re_inst_2_io_op1; // @[Float.scala 45:22]
  wire [16:0] io_res_re_inst_2_io_op2; // @[Float.scala 45:22]
  wire [16:0] io_res_re_inst_2_io_res; // @[Float.scala 45:22]
  wire [16:0] io_res_im_inst_io_op1; // @[Float.scala 64:22]
  wire [16:0] io_res_im_inst_io_op2; // @[Float.scala 64:22]
  wire [16:0] io_res_im_inst_io_res; // @[Float.scala 64:22]
  wire [16:0] io_res_im_inst_1_io_op1; // @[Float.scala 64:22]
  wire [16:0] io_res_im_inst_1_io_op2; // @[Float.scala 64:22]
  wire [16:0] io_res_im_inst_1_io_res; // @[Float.scala 64:22]
  wire [16:0] io_res_im_inst_2_io_op1; // @[Float.scala 25:22]
  wire [16:0] io_res_im_inst_2_io_op2; // @[Float.scala 25:22]
  wire [16:0] io_res_im_inst_2_io_res; // @[Float.scala 25:22]
  FloatMul io_res_re_inst ( // @[Float.scala 64:22]
    .io_op1(io_res_re_inst_io_op1),
    .io_op2(io_res_re_inst_io_op2),
    .io_res(io_res_re_inst_io_res)
  );
  FloatMul io_res_re_inst_1 ( // @[Float.scala 64:22]
    .io_op1(io_res_re_inst_1_io_op1),
    .io_op2(io_res_re_inst_1_io_op2),
    .io_res(io_res_re_inst_1_io_res)
  );
  FloatSub io_res_re_inst_2 ( // @[Float.scala 45:22]
    .io_op1(io_res_re_inst_2_io_op1),
    .io_op2(io_res_re_inst_2_io_op2),
    .io_res(io_res_re_inst_2_io_res)
  );
  FloatMul io_res_im_inst ( // @[Float.scala 64:22]
    .io_op1(io_res_im_inst_io_op1),
    .io_op2(io_res_im_inst_io_op2),
    .io_res(io_res_im_inst_io_res)
  );
  FloatMul io_res_im_inst_1 ( // @[Float.scala 64:22]
    .io_op1(io_res_im_inst_1_io_op1),
    .io_op2(io_res_im_inst_1_io_op2),
    .io_res(io_res_im_inst_1_io_res)
  );
  FloatAdd io_res_im_inst_2 ( // @[Float.scala 25:22]
    .io_op1(io_res_im_inst_2_io_op1),
    .io_op2(io_res_im_inst_2_io_op2),
    .io_res(io_res_im_inst_2_io_res)
  );
  assign io_res_re = io_res_re_inst_2_io_res; // @[Modules.scala 139:17]
  assign io_res_im = io_res_im_inst_2_io_res; // @[Modules.scala 140:17]
  assign io_res_re_inst_io_op1 = io_op1_re; // @[Float.scala 65:17]
  assign io_res_re_inst_io_op2 = io_op2_re; // @[Float.scala 66:17]
  assign io_res_re_inst_1_io_op1 = io_op1_im; // @[Float.scala 65:17]
  assign io_res_re_inst_1_io_op2 = io_op2_im; // @[Float.scala 66:17]
  assign io_res_re_inst_2_io_op1 = io_res_re_inst_io_res; // @[Float.scala 46:17]
  assign io_res_re_inst_2_io_op2 = io_res_re_inst_1_io_res; // @[Float.scala 47:17]
  assign io_res_im_inst_io_op1 = io_op1_re; // @[Float.scala 65:17]
  assign io_res_im_inst_io_op2 = io_op2_im; // @[Float.scala 66:17]
  assign io_res_im_inst_1_io_op1 = io_op1_im; // @[Float.scala 65:17]
  assign io_res_im_inst_1_io_op2 = io_op2_re; // @[Float.scala 66:17]
  assign io_res_im_inst_2_io_op1 = io_res_im_inst_io_res; // @[Float.scala 26:17]
  assign io_res_im_inst_2_io_op2 = io_res_im_inst_1_io_res; // @[Float.scala 27:17]
endmodule
module ButterflyMul(
  input  [16:0] io_in_0_re,
  input  [16:0] io_in_0_im,
  input  [16:0] io_in_1_re,
  input  [16:0] io_in_1_im,
  output [16:0] io_out_0_re,
  output [16:0] io_out_0_im,
  output [16:0] io_out_1_re,
  output [16:0] io_out_1_im,
  input  [16:0] io_wn_0_re,
  input  [16:0] io_wn_0_im
);
  wire [16:0] temp_0_inst_io_op1_re; // @[Modules.scala 81:22]
  wire [16:0] temp_0_inst_io_op1_im; // @[Modules.scala 81:22]
  wire [16:0] temp_0_inst_io_op2_re; // @[Modules.scala 81:22]
  wire [16:0] temp_0_inst_io_op2_im; // @[Modules.scala 81:22]
  wire [16:0] temp_0_inst_io_res_re; // @[Modules.scala 81:22]
  wire [16:0] temp_0_inst_io_res_im; // @[Modules.scala 81:22]
  wire [16:0] temp_1_inst_io_op1_re; // @[Modules.scala 100:22]
  wire [16:0] temp_1_inst_io_op1_im; // @[Modules.scala 100:22]
  wire [16:0] temp_1_inst_io_op2_re; // @[Modules.scala 100:22]
  wire [16:0] temp_1_inst_io_op2_im; // @[Modules.scala 100:22]
  wire [16:0] temp_1_inst_io_res_re; // @[Modules.scala 100:22]
  wire [16:0] temp_1_inst_io_res_im; // @[Modules.scala 100:22]
  wire [16:0] io_out_1_inst_io_op1_re; // @[Modules.scala 158:22]
  wire [16:0] io_out_1_inst_io_op1_im; // @[Modules.scala 158:22]
  wire [16:0] io_out_1_inst_io_op2_re; // @[Modules.scala 158:22]
  wire [16:0] io_out_1_inst_io_op2_im; // @[Modules.scala 158:22]
  wire [16:0] io_out_1_inst_io_res_re; // @[Modules.scala 158:22]
  wire [16:0] io_out_1_inst_io_res_im; // @[Modules.scala 158:22]
  ComplexAdd temp_0_inst ( // @[Modules.scala 81:22]
    .io_op1_re(temp_0_inst_io_op1_re),
    .io_op1_im(temp_0_inst_io_op1_im),
    .io_op2_re(temp_0_inst_io_op2_re),
    .io_op2_im(temp_0_inst_io_op2_im),
    .io_res_re(temp_0_inst_io_res_re),
    .io_res_im(temp_0_inst_io_res_im)
  );
  ComplexSub temp_1_inst ( // @[Modules.scala 100:22]
    .io_op1_re(temp_1_inst_io_op1_re),
    .io_op1_im(temp_1_inst_io_op1_im),
    .io_op2_re(temp_1_inst_io_op2_re),
    .io_op2_im(temp_1_inst_io_op2_im),
    .io_res_re(temp_1_inst_io_res_re),
    .io_res_im(temp_1_inst_io_res_im)
  );
  ComplexMul io_out_1_inst ( // @[Modules.scala 158:22]
    .io_op1_re(io_out_1_inst_io_op1_re),
    .io_op1_im(io_out_1_inst_io_op1_im),
    .io_op2_re(io_out_1_inst_io_op2_re),
    .io_op2_im(io_out_1_inst_io_op2_im),
    .io_res_re(io_out_1_inst_io_res_re),
    .io_res_im(io_out_1_inst_io_res_im)
  );
  assign io_out_0_re = temp_0_inst_io_res_re; // @[Modules.scala 224:21 226:13]
  assign io_out_0_im = temp_0_inst_io_res_im; // @[Modules.scala 224:21 226:13]
  assign io_out_1_re = io_out_1_inst_io_res_re; // @[Modules.scala 267:15]
  assign io_out_1_im = io_out_1_inst_io_res_im; // @[Modules.scala 267:15]
  assign temp_0_inst_io_op1_re = io_in_0_re; // @[Modules.scala 82:17]
  assign temp_0_inst_io_op1_im = io_in_0_im; // @[Modules.scala 82:17]
  assign temp_0_inst_io_op2_re = io_in_1_re; // @[Modules.scala 83:17]
  assign temp_0_inst_io_op2_im = io_in_1_im; // @[Modules.scala 83:17]
  assign temp_1_inst_io_op1_re = io_in_0_re; // @[Modules.scala 101:17]
  assign temp_1_inst_io_op1_im = io_in_0_im; // @[Modules.scala 101:17]
  assign temp_1_inst_io_op2_re = io_in_1_re; // @[Modules.scala 102:17]
  assign temp_1_inst_io_op2_im = io_in_1_im; // @[Modules.scala 102:17]
  assign io_out_1_inst_io_op1_re = temp_1_inst_io_res_re; // @[Modules.scala 224:21 227:13]
  assign io_out_1_inst_io_op1_im = temp_1_inst_io_res_im; // @[Modules.scala 224:21 227:13]
  assign io_out_1_inst_io_op2_re = io_wn_0_re; // @[Modules.scala 160:17]
  assign io_out_1_inst_io_op2_im = io_wn_0_im; // @[Modules.scala 160:17]
endmodule
module ButterflyAdd(
  input  [16:0] io_in_0_re,
  input  [16:0] io_in_0_im,
  input  [16:0] io_in_1_re,
  input  [16:0] io_in_1_im,
  output [16:0] io_out_0_re,
  output [16:0] io_out_0_im,
  output [16:0] io_out_1_re,
  output [16:0] io_out_1_im
);
  wire [16:0] io_out_0_inst_io_op1_re; // @[Modules.scala 81:22]
  wire [16:0] io_out_0_inst_io_op1_im; // @[Modules.scala 81:22]
  wire [16:0] io_out_0_inst_io_op2_re; // @[Modules.scala 81:22]
  wire [16:0] io_out_0_inst_io_op2_im; // @[Modules.scala 81:22]
  wire [16:0] io_out_0_inst_io_res_re; // @[Modules.scala 81:22]
  wire [16:0] io_out_0_inst_io_res_im; // @[Modules.scala 81:22]
  wire [16:0] io_out_1_inst_io_op1_re; // @[Modules.scala 100:22]
  wire [16:0] io_out_1_inst_io_op1_im; // @[Modules.scala 100:22]
  wire [16:0] io_out_1_inst_io_op2_re; // @[Modules.scala 100:22]
  wire [16:0] io_out_1_inst_io_op2_im; // @[Modules.scala 100:22]
  wire [16:0] io_out_1_inst_io_res_re; // @[Modules.scala 100:22]
  wire [16:0] io_out_1_inst_io_res_im; // @[Modules.scala 100:22]
  ComplexAdd io_out_0_inst ( // @[Modules.scala 81:22]
    .io_op1_re(io_out_0_inst_io_op1_re),
    .io_op1_im(io_out_0_inst_io_op1_im),
    .io_op2_re(io_out_0_inst_io_op2_re),
    .io_op2_im(io_out_0_inst_io_op2_im),
    .io_res_re(io_out_0_inst_io_res_re),
    .io_res_im(io_out_0_inst_io_res_im)
  );
  ComplexSub io_out_1_inst ( // @[Modules.scala 100:22]
    .io_op1_re(io_out_1_inst_io_op1_re),
    .io_op1_im(io_out_1_inst_io_op1_im),
    .io_op2_re(io_out_1_inst_io_op2_re),
    .io_op2_im(io_out_1_inst_io_op2_im),
    .io_res_re(io_out_1_inst_io_res_re),
    .io_res_im(io_out_1_inst_io_res_im)
  );
  assign io_out_0_re = io_out_0_inst_io_res_re; // @[Modules.scala 170:15]
  assign io_out_0_im = io_out_0_inst_io_res_im; // @[Modules.scala 170:15]
  assign io_out_1_re = io_out_1_inst_io_res_re; // @[Modules.scala 171:15]
  assign io_out_1_im = io_out_1_inst_io_res_im; // @[Modules.scala 171:15]
  assign io_out_0_inst_io_op1_re = io_in_0_re; // @[Modules.scala 82:17]
  assign io_out_0_inst_io_op1_im = io_in_0_im; // @[Modules.scala 82:17]
  assign io_out_0_inst_io_op2_re = io_in_1_re; // @[Modules.scala 83:17]
  assign io_out_0_inst_io_op2_im = io_in_1_im; // @[Modules.scala 83:17]
  assign io_out_1_inst_io_op1_re = io_in_0_re; // @[Modules.scala 101:17]
  assign io_out_1_inst_io_op1_im = io_in_0_im; // @[Modules.scala 101:17]
  assign io_out_1_inst_io_op2_re = io_in_1_re; // @[Modules.scala 102:17]
  assign io_out_1_inst_io_op2_im = io_in_1_im; // @[Modules.scala 102:17]
endmodule
module Switch(
  input         clock,
  input  [16:0] io_in_0_re,
  input  [16:0] io_in_0_im,
  input  [16:0] io_in_1_re,
  input  [16:0] io_in_1_im,
  output [16:0] io_out_0_re,
  output [16:0] io_out_0_im,
  output [16:0] io_out_1_re,
  output [16:0] io_out_1_im,
  input         io_sel
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_9;
  reg [31:0] _RAND_10;
  reg [31:0] _RAND_11;
  reg [31:0] _RAND_12;
  reg [31:0] _RAND_13;
  reg [31:0] _RAND_14;
  reg [31:0] _RAND_15;
  reg [31:0] _RAND_16;
  reg [31:0] _RAND_17;
  reg [31:0] _RAND_18;
  reg [31:0] _RAND_19;
  reg [31:0] _RAND_20;
  reg [31:0] _RAND_21;
  reg [31:0] _RAND_22;
  reg [31:0] _RAND_23;
  reg [31:0] _RAND_24;
  reg [31:0] _RAND_25;
  reg [31:0] _RAND_26;
  reg [31:0] _RAND_27;
  reg [31:0] _RAND_28;
  reg [31:0] _RAND_29;
  reg [31:0] _RAND_30;
  reg [31:0] _RAND_31;
  reg [31:0] _RAND_32;
  reg [31:0] _RAND_33;
  reg [31:0] _RAND_34;
  reg [31:0] _RAND_35;
  reg [31:0] _RAND_36;
  reg [31:0] _RAND_37;
  reg [31:0] _RAND_38;
  reg [31:0] _RAND_39;
  reg [31:0] _RAND_40;
  reg [31:0] _RAND_41;
  reg [31:0] _RAND_42;
  reg [31:0] _RAND_43;
  reg [31:0] _RAND_44;
  reg [31:0] _RAND_45;
  reg [31:0] _RAND_46;
  reg [31:0] _RAND_47;
  reg [31:0] _RAND_48;
  reg [31:0] _RAND_49;
  reg [31:0] _RAND_50;
  reg [31:0] _RAND_51;
  reg [31:0] _RAND_52;
  reg [31:0] _RAND_53;
  reg [31:0] _RAND_54;
  reg [31:0] _RAND_55;
  reg [31:0] _RAND_56;
  reg [31:0] _RAND_57;
  reg [31:0] _RAND_58;
  reg [31:0] _RAND_59;
  reg [31:0] _RAND_60;
  reg [31:0] _RAND_61;
  reg [31:0] _RAND_62;
  reg [31:0] _RAND_63;
  reg [31:0] _RAND_64;
  reg [31:0] _RAND_65;
  reg [31:0] _RAND_66;
  reg [31:0] _RAND_67;
  reg [31:0] _RAND_68;
  reg [31:0] _RAND_69;
  reg [31:0] _RAND_70;
  reg [31:0] _RAND_71;
  reg [31:0] _RAND_72;
  reg [31:0] _RAND_73;
  reg [31:0] _RAND_74;
  reg [31:0] _RAND_75;
  reg [31:0] _RAND_76;
  reg [31:0] _RAND_77;
  reg [31:0] _RAND_78;
  reg [31:0] _RAND_79;
  reg [31:0] _RAND_80;
  reg [31:0] _RAND_81;
  reg [31:0] _RAND_82;
  reg [31:0] _RAND_83;
  reg [31:0] _RAND_84;
  reg [31:0] _RAND_85;
  reg [31:0] _RAND_86;
  reg [31:0] _RAND_87;
  reg [31:0] _RAND_88;
  reg [31:0] _RAND_89;
  reg [31:0] _RAND_90;
  reg [31:0] _RAND_91;
  reg [31:0] _RAND_92;
  reg [31:0] _RAND_93;
  reg [31:0] _RAND_94;
  reg [31:0] _RAND_95;
  reg [31:0] _RAND_96;
  reg [31:0] _RAND_97;
  reg [31:0] _RAND_98;
  reg [31:0] _RAND_99;
  reg [31:0] _RAND_100;
  reg [31:0] _RAND_101;
  reg [31:0] _RAND_102;
  reg [31:0] _RAND_103;
  reg [31:0] _RAND_104;
  reg [31:0] _RAND_105;
  reg [31:0] _RAND_106;
  reg [31:0] _RAND_107;
  reg [31:0] _RAND_108;
  reg [31:0] _RAND_109;
  reg [31:0] _RAND_110;
  reg [31:0] _RAND_111;
  reg [31:0] _RAND_112;
  reg [31:0] _RAND_113;
  reg [31:0] _RAND_114;
  reg [31:0] _RAND_115;
  reg [31:0] _RAND_116;
  reg [31:0] _RAND_117;
  reg [31:0] _RAND_118;
  reg [31:0] _RAND_119;
  reg [31:0] _RAND_120;
  reg [31:0] _RAND_121;
  reg [31:0] _RAND_122;
  reg [31:0] _RAND_123;
  reg [31:0] _RAND_124;
  reg [31:0] _RAND_125;
  reg [31:0] _RAND_126;
  reg [31:0] _RAND_127;
  reg [31:0] _RAND_128;
  reg [31:0] _RAND_129;
  reg [31:0] _RAND_130;
  reg [31:0] _RAND_131;
  reg [31:0] _RAND_132;
  reg [31:0] _RAND_133;
  reg [31:0] _RAND_134;
  reg [31:0] _RAND_135;
  reg [31:0] _RAND_136;
  reg [31:0] _RAND_137;
  reg [31:0] _RAND_138;
  reg [31:0] _RAND_139;
  reg [31:0] _RAND_140;
  reg [31:0] _RAND_141;
  reg [31:0] _RAND_142;
  reg [31:0] _RAND_143;
  reg [31:0] _RAND_144;
  reg [31:0] _RAND_145;
  reg [31:0] _RAND_146;
  reg [31:0] _RAND_147;
  reg [31:0] _RAND_148;
  reg [31:0] _RAND_149;
  reg [31:0] _RAND_150;
  reg [31:0] _RAND_151;
  reg [31:0] _RAND_152;
  reg [31:0] _RAND_153;
  reg [31:0] _RAND_154;
  reg [31:0] _RAND_155;
  reg [31:0] _RAND_156;
  reg [31:0] _RAND_157;
  reg [31:0] _RAND_158;
  reg [31:0] _RAND_159;
  reg [31:0] _RAND_160;
  reg [31:0] _RAND_161;
  reg [31:0] _RAND_162;
  reg [31:0] _RAND_163;
  reg [31:0] _RAND_164;
  reg [31:0] _RAND_165;
  reg [31:0] _RAND_166;
  reg [31:0] _RAND_167;
  reg [31:0] _RAND_168;
  reg [31:0] _RAND_169;
  reg [31:0] _RAND_170;
  reg [31:0] _RAND_171;
  reg [31:0] _RAND_172;
  reg [31:0] _RAND_173;
  reg [31:0] _RAND_174;
  reg [31:0] _RAND_175;
  reg [31:0] _RAND_176;
  reg [31:0] _RAND_177;
  reg [31:0] _RAND_178;
  reg [31:0] _RAND_179;
  reg [31:0] _RAND_180;
  reg [31:0] _RAND_181;
  reg [31:0] _RAND_182;
  reg [31:0] _RAND_183;
  reg [31:0] _RAND_184;
  reg [31:0] _RAND_185;
  reg [31:0] _RAND_186;
  reg [31:0] _RAND_187;
  reg [31:0] _RAND_188;
  reg [31:0] _RAND_189;
  reg [31:0] _RAND_190;
  reg [31:0] _RAND_191;
  reg [31:0] _RAND_192;
  reg [31:0] _RAND_193;
  reg [31:0] _RAND_194;
  reg [31:0] _RAND_195;
  reg [31:0] _RAND_196;
  reg [31:0] _RAND_197;
  reg [31:0] _RAND_198;
  reg [31:0] _RAND_199;
  reg [31:0] _RAND_200;
  reg [31:0] _RAND_201;
  reg [31:0] _RAND_202;
  reg [31:0] _RAND_203;
  reg [31:0] _RAND_204;
  reg [31:0] _RAND_205;
  reg [31:0] _RAND_206;
  reg [31:0] _RAND_207;
  reg [31:0] _RAND_208;
  reg [31:0] _RAND_209;
  reg [31:0] _RAND_210;
  reg [31:0] _RAND_211;
  reg [31:0] _RAND_212;
  reg [31:0] _RAND_213;
  reg [31:0] _RAND_214;
  reg [31:0] _RAND_215;
  reg [31:0] _RAND_216;
  reg [31:0] _RAND_217;
  reg [31:0] _RAND_218;
  reg [31:0] _RAND_219;
  reg [31:0] _RAND_220;
  reg [31:0] _RAND_221;
  reg [31:0] _RAND_222;
  reg [31:0] _RAND_223;
  reg [31:0] _RAND_224;
  reg [31:0] _RAND_225;
  reg [31:0] _RAND_226;
  reg [31:0] _RAND_227;
  reg [31:0] _RAND_228;
  reg [31:0] _RAND_229;
  reg [31:0] _RAND_230;
  reg [31:0] _RAND_231;
  reg [31:0] _RAND_232;
  reg [31:0] _RAND_233;
  reg [31:0] _RAND_234;
  reg [31:0] _RAND_235;
  reg [31:0] _RAND_236;
  reg [31:0] _RAND_237;
  reg [31:0] _RAND_238;
  reg [31:0] _RAND_239;
  reg [31:0] _RAND_240;
  reg [31:0] _RAND_241;
  reg [31:0] _RAND_242;
  reg [31:0] _RAND_243;
  reg [31:0] _RAND_244;
  reg [31:0] _RAND_245;
  reg [31:0] _RAND_246;
  reg [31:0] _RAND_247;
  reg [31:0] _RAND_248;
  reg [31:0] _RAND_249;
  reg [31:0] _RAND_250;
  reg [31:0] _RAND_251;
  reg [31:0] _RAND_252;
  reg [31:0] _RAND_253;
  reg [31:0] _RAND_254;
  reg [31:0] _RAND_255;
`endif // RANDOMIZE_REG_INIT
  reg [16:0] swdata_1_r_re; // @[Reg.scala 19:16]
  reg [16:0] swdata_1_r_im; // @[Reg.scala 19:16]
  reg [16:0] swdata_1_r_1_re; // @[Reg.scala 19:16]
  reg [16:0] swdata_1_r_1_im; // @[Reg.scala 19:16]
  reg [16:0] swdata_1_r_2_re; // @[Reg.scala 19:16]
  reg [16:0] swdata_1_r_2_im; // @[Reg.scala 19:16]
  reg [16:0] swdata_1_r_3_re; // @[Reg.scala 19:16]
  reg [16:0] swdata_1_r_3_im; // @[Reg.scala 19:16]
  reg [16:0] swdata_1_r_4_re; // @[Reg.scala 19:16]
  reg [16:0] swdata_1_r_4_im; // @[Reg.scala 19:16]
  reg [16:0] swdata_1_r_5_re; // @[Reg.scala 19:16]
  reg [16:0] swdata_1_r_5_im; // @[Reg.scala 19:16]
  reg [16:0] swdata_1_r_6_re; // @[Reg.scala 19:16]
  reg [16:0] swdata_1_r_6_im; // @[Reg.scala 19:16]
  reg [16:0] swdata_1_r_7_re; // @[Reg.scala 19:16]
  reg [16:0] swdata_1_r_7_im; // @[Reg.scala 19:16]
  reg [16:0] swdata_1_r_8_re; // @[Reg.scala 19:16]
  reg [16:0] swdata_1_r_8_im; // @[Reg.scala 19:16]
  reg [16:0] swdata_1_r_9_re; // @[Reg.scala 19:16]
  reg [16:0] swdata_1_r_9_im; // @[Reg.scala 19:16]
  reg [16:0] swdata_1_r_10_re; // @[Reg.scala 19:16]
  reg [16:0] swdata_1_r_10_im; // @[Reg.scala 19:16]
  reg [16:0] swdata_1_r_11_re; // @[Reg.scala 19:16]
  reg [16:0] swdata_1_r_11_im; // @[Reg.scala 19:16]
  reg [16:0] swdata_1_r_12_re; // @[Reg.scala 19:16]
  reg [16:0] swdata_1_r_12_im; // @[Reg.scala 19:16]
  reg [16:0] swdata_1_r_13_re; // @[Reg.scala 19:16]
  reg [16:0] swdata_1_r_13_im; // @[Reg.scala 19:16]
  reg [16:0] swdata_1_r_14_re; // @[Reg.scala 19:16]
  reg [16:0] swdata_1_r_14_im; // @[Reg.scala 19:16]
  reg [16:0] swdata_1_r_15_re; // @[Reg.scala 19:16]
  reg [16:0] swdata_1_r_15_im; // @[Reg.scala 19:16]
  reg [16:0] swdata_1_r_16_re; // @[Reg.scala 19:16]
  reg [16:0] swdata_1_r_16_im; // @[Reg.scala 19:16]
  reg [16:0] swdata_1_r_17_re; // @[Reg.scala 19:16]
  reg [16:0] swdata_1_r_17_im; // @[Reg.scala 19:16]
  reg [16:0] swdata_1_r_18_re; // @[Reg.scala 19:16]
  reg [16:0] swdata_1_r_18_im; // @[Reg.scala 19:16]
  reg [16:0] swdata_1_r_19_re; // @[Reg.scala 19:16]
  reg [16:0] swdata_1_r_19_im; // @[Reg.scala 19:16]
  reg [16:0] swdata_1_r_20_re; // @[Reg.scala 19:16]
  reg [16:0] swdata_1_r_20_im; // @[Reg.scala 19:16]
  reg [16:0] swdata_1_r_21_re; // @[Reg.scala 19:16]
  reg [16:0] swdata_1_r_21_im; // @[Reg.scala 19:16]
  reg [16:0] swdata_1_r_22_re; // @[Reg.scala 19:16]
  reg [16:0] swdata_1_r_22_im; // @[Reg.scala 19:16]
  reg [16:0] swdata_1_r_23_re; // @[Reg.scala 19:16]
  reg [16:0] swdata_1_r_23_im; // @[Reg.scala 19:16]
  reg [16:0] swdata_1_r_24_re; // @[Reg.scala 19:16]
  reg [16:0] swdata_1_r_24_im; // @[Reg.scala 19:16]
  reg [16:0] swdata_1_r_25_re; // @[Reg.scala 19:16]
  reg [16:0] swdata_1_r_25_im; // @[Reg.scala 19:16]
  reg [16:0] swdata_1_r_26_re; // @[Reg.scala 19:16]
  reg [16:0] swdata_1_r_26_im; // @[Reg.scala 19:16]
  reg [16:0] swdata_1_r_27_re; // @[Reg.scala 19:16]
  reg [16:0] swdata_1_r_27_im; // @[Reg.scala 19:16]
  reg [16:0] swdata_1_r_28_re; // @[Reg.scala 19:16]
  reg [16:0] swdata_1_r_28_im; // @[Reg.scala 19:16]
  reg [16:0] swdata_1_r_29_re; // @[Reg.scala 19:16]
  reg [16:0] swdata_1_r_29_im; // @[Reg.scala 19:16]
  reg [16:0] swdata_1_r_30_re; // @[Reg.scala 19:16]
  reg [16:0] swdata_1_r_30_im; // @[Reg.scala 19:16]
  reg [16:0] swdata_1_r_31_re; // @[Reg.scala 19:16]
  reg [16:0] swdata_1_r_31_im; // @[Reg.scala 19:16]
  reg [16:0] swdata_1_r_32_re; // @[Reg.scala 19:16]
  reg [16:0] swdata_1_r_32_im; // @[Reg.scala 19:16]
  reg [16:0] swdata_1_r_33_re; // @[Reg.scala 19:16]
  reg [16:0] swdata_1_r_33_im; // @[Reg.scala 19:16]
  reg [16:0] swdata_1_r_34_re; // @[Reg.scala 19:16]
  reg [16:0] swdata_1_r_34_im; // @[Reg.scala 19:16]
  reg [16:0] swdata_1_r_35_re; // @[Reg.scala 19:16]
  reg [16:0] swdata_1_r_35_im; // @[Reg.scala 19:16]
  reg [16:0] swdata_1_r_36_re; // @[Reg.scala 19:16]
  reg [16:0] swdata_1_r_36_im; // @[Reg.scala 19:16]
  reg [16:0] swdata_1_r_37_re; // @[Reg.scala 19:16]
  reg [16:0] swdata_1_r_37_im; // @[Reg.scala 19:16]
  reg [16:0] swdata_1_r_38_re; // @[Reg.scala 19:16]
  reg [16:0] swdata_1_r_38_im; // @[Reg.scala 19:16]
  reg [16:0] swdata_1_r_39_re; // @[Reg.scala 19:16]
  reg [16:0] swdata_1_r_39_im; // @[Reg.scala 19:16]
  reg [16:0] swdata_1_r_40_re; // @[Reg.scala 19:16]
  reg [16:0] swdata_1_r_40_im; // @[Reg.scala 19:16]
  reg [16:0] swdata_1_r_41_re; // @[Reg.scala 19:16]
  reg [16:0] swdata_1_r_41_im; // @[Reg.scala 19:16]
  reg [16:0] swdata_1_r_42_re; // @[Reg.scala 19:16]
  reg [16:0] swdata_1_r_42_im; // @[Reg.scala 19:16]
  reg [16:0] swdata_1_r_43_re; // @[Reg.scala 19:16]
  reg [16:0] swdata_1_r_43_im; // @[Reg.scala 19:16]
  reg [16:0] swdata_1_r_44_re; // @[Reg.scala 19:16]
  reg [16:0] swdata_1_r_44_im; // @[Reg.scala 19:16]
  reg [16:0] swdata_1_r_45_re; // @[Reg.scala 19:16]
  reg [16:0] swdata_1_r_45_im; // @[Reg.scala 19:16]
  reg [16:0] swdata_1_r_46_re; // @[Reg.scala 19:16]
  reg [16:0] swdata_1_r_46_im; // @[Reg.scala 19:16]
  reg [16:0] swdata_1_r_47_re; // @[Reg.scala 19:16]
  reg [16:0] swdata_1_r_47_im; // @[Reg.scala 19:16]
  reg [16:0] swdata_1_r_48_re; // @[Reg.scala 19:16]
  reg [16:0] swdata_1_r_48_im; // @[Reg.scala 19:16]
  reg [16:0] swdata_1_r_49_re; // @[Reg.scala 19:16]
  reg [16:0] swdata_1_r_49_im; // @[Reg.scala 19:16]
  reg [16:0] swdata_1_r_50_re; // @[Reg.scala 19:16]
  reg [16:0] swdata_1_r_50_im; // @[Reg.scala 19:16]
  reg [16:0] swdata_1_r_51_re; // @[Reg.scala 19:16]
  reg [16:0] swdata_1_r_51_im; // @[Reg.scala 19:16]
  reg [16:0] swdata_1_r_52_re; // @[Reg.scala 19:16]
  reg [16:0] swdata_1_r_52_im; // @[Reg.scala 19:16]
  reg [16:0] swdata_1_r_53_re; // @[Reg.scala 19:16]
  reg [16:0] swdata_1_r_53_im; // @[Reg.scala 19:16]
  reg [16:0] swdata_1_r_54_re; // @[Reg.scala 19:16]
  reg [16:0] swdata_1_r_54_im; // @[Reg.scala 19:16]
  reg [16:0] swdata_1_r_55_re; // @[Reg.scala 19:16]
  reg [16:0] swdata_1_r_55_im; // @[Reg.scala 19:16]
  reg [16:0] swdata_1_r_56_re; // @[Reg.scala 19:16]
  reg [16:0] swdata_1_r_56_im; // @[Reg.scala 19:16]
  reg [16:0] swdata_1_r_57_re; // @[Reg.scala 19:16]
  reg [16:0] swdata_1_r_57_im; // @[Reg.scala 19:16]
  reg [16:0] swdata_1_r_58_re; // @[Reg.scala 19:16]
  reg [16:0] swdata_1_r_58_im; // @[Reg.scala 19:16]
  reg [16:0] swdata_1_r_59_re; // @[Reg.scala 19:16]
  reg [16:0] swdata_1_r_59_im; // @[Reg.scala 19:16]
  reg [16:0] swdata_1_r_60_re; // @[Reg.scala 19:16]
  reg [16:0] swdata_1_r_60_im; // @[Reg.scala 19:16]
  reg [16:0] swdata_1_r_61_re; // @[Reg.scala 19:16]
  reg [16:0] swdata_1_r_61_im; // @[Reg.scala 19:16]
  reg [16:0] swdata_1_r_62_re; // @[Reg.scala 19:16]
  reg [16:0] swdata_1_r_62_im; // @[Reg.scala 19:16]
  reg [16:0] swdata_1_r_63_re; // @[Reg.scala 19:16]
  reg [16:0] swdata_1_r_63_im; // @[Reg.scala 19:16]
  reg [16:0] io_out_0_r_re; // @[Reg.scala 19:16]
  reg [16:0] io_out_0_r_im; // @[Reg.scala 19:16]
  reg [16:0] io_out_0_r_1_re; // @[Reg.scala 19:16]
  reg [16:0] io_out_0_r_1_im; // @[Reg.scala 19:16]
  reg [16:0] io_out_0_r_2_re; // @[Reg.scala 19:16]
  reg [16:0] io_out_0_r_2_im; // @[Reg.scala 19:16]
  reg [16:0] io_out_0_r_3_re; // @[Reg.scala 19:16]
  reg [16:0] io_out_0_r_3_im; // @[Reg.scala 19:16]
  reg [16:0] io_out_0_r_4_re; // @[Reg.scala 19:16]
  reg [16:0] io_out_0_r_4_im; // @[Reg.scala 19:16]
  reg [16:0] io_out_0_r_5_re; // @[Reg.scala 19:16]
  reg [16:0] io_out_0_r_5_im; // @[Reg.scala 19:16]
  reg [16:0] io_out_0_r_6_re; // @[Reg.scala 19:16]
  reg [16:0] io_out_0_r_6_im; // @[Reg.scala 19:16]
  reg [16:0] io_out_0_r_7_re; // @[Reg.scala 19:16]
  reg [16:0] io_out_0_r_7_im; // @[Reg.scala 19:16]
  reg [16:0] io_out_0_r_8_re; // @[Reg.scala 19:16]
  reg [16:0] io_out_0_r_8_im; // @[Reg.scala 19:16]
  reg [16:0] io_out_0_r_9_re; // @[Reg.scala 19:16]
  reg [16:0] io_out_0_r_9_im; // @[Reg.scala 19:16]
  reg [16:0] io_out_0_r_10_re; // @[Reg.scala 19:16]
  reg [16:0] io_out_0_r_10_im; // @[Reg.scala 19:16]
  reg [16:0] io_out_0_r_11_re; // @[Reg.scala 19:16]
  reg [16:0] io_out_0_r_11_im; // @[Reg.scala 19:16]
  reg [16:0] io_out_0_r_12_re; // @[Reg.scala 19:16]
  reg [16:0] io_out_0_r_12_im; // @[Reg.scala 19:16]
  reg [16:0] io_out_0_r_13_re; // @[Reg.scala 19:16]
  reg [16:0] io_out_0_r_13_im; // @[Reg.scala 19:16]
  reg [16:0] io_out_0_r_14_re; // @[Reg.scala 19:16]
  reg [16:0] io_out_0_r_14_im; // @[Reg.scala 19:16]
  reg [16:0] io_out_0_r_15_re; // @[Reg.scala 19:16]
  reg [16:0] io_out_0_r_15_im; // @[Reg.scala 19:16]
  reg [16:0] io_out_0_r_16_re; // @[Reg.scala 19:16]
  reg [16:0] io_out_0_r_16_im; // @[Reg.scala 19:16]
  reg [16:0] io_out_0_r_17_re; // @[Reg.scala 19:16]
  reg [16:0] io_out_0_r_17_im; // @[Reg.scala 19:16]
  reg [16:0] io_out_0_r_18_re; // @[Reg.scala 19:16]
  reg [16:0] io_out_0_r_18_im; // @[Reg.scala 19:16]
  reg [16:0] io_out_0_r_19_re; // @[Reg.scala 19:16]
  reg [16:0] io_out_0_r_19_im; // @[Reg.scala 19:16]
  reg [16:0] io_out_0_r_20_re; // @[Reg.scala 19:16]
  reg [16:0] io_out_0_r_20_im; // @[Reg.scala 19:16]
  reg [16:0] io_out_0_r_21_re; // @[Reg.scala 19:16]
  reg [16:0] io_out_0_r_21_im; // @[Reg.scala 19:16]
  reg [16:0] io_out_0_r_22_re; // @[Reg.scala 19:16]
  reg [16:0] io_out_0_r_22_im; // @[Reg.scala 19:16]
  reg [16:0] io_out_0_r_23_re; // @[Reg.scala 19:16]
  reg [16:0] io_out_0_r_23_im; // @[Reg.scala 19:16]
  reg [16:0] io_out_0_r_24_re; // @[Reg.scala 19:16]
  reg [16:0] io_out_0_r_24_im; // @[Reg.scala 19:16]
  reg [16:0] io_out_0_r_25_re; // @[Reg.scala 19:16]
  reg [16:0] io_out_0_r_25_im; // @[Reg.scala 19:16]
  reg [16:0] io_out_0_r_26_re; // @[Reg.scala 19:16]
  reg [16:0] io_out_0_r_26_im; // @[Reg.scala 19:16]
  reg [16:0] io_out_0_r_27_re; // @[Reg.scala 19:16]
  reg [16:0] io_out_0_r_27_im; // @[Reg.scala 19:16]
  reg [16:0] io_out_0_r_28_re; // @[Reg.scala 19:16]
  reg [16:0] io_out_0_r_28_im; // @[Reg.scala 19:16]
  reg [16:0] io_out_0_r_29_re; // @[Reg.scala 19:16]
  reg [16:0] io_out_0_r_29_im; // @[Reg.scala 19:16]
  reg [16:0] io_out_0_r_30_re; // @[Reg.scala 19:16]
  reg [16:0] io_out_0_r_30_im; // @[Reg.scala 19:16]
  reg [16:0] io_out_0_r_31_re; // @[Reg.scala 19:16]
  reg [16:0] io_out_0_r_31_im; // @[Reg.scala 19:16]
  reg [16:0] io_out_0_r_32_re; // @[Reg.scala 19:16]
  reg [16:0] io_out_0_r_32_im; // @[Reg.scala 19:16]
  reg [16:0] io_out_0_r_33_re; // @[Reg.scala 19:16]
  reg [16:0] io_out_0_r_33_im; // @[Reg.scala 19:16]
  reg [16:0] io_out_0_r_34_re; // @[Reg.scala 19:16]
  reg [16:0] io_out_0_r_34_im; // @[Reg.scala 19:16]
  reg [16:0] io_out_0_r_35_re; // @[Reg.scala 19:16]
  reg [16:0] io_out_0_r_35_im; // @[Reg.scala 19:16]
  reg [16:0] io_out_0_r_36_re; // @[Reg.scala 19:16]
  reg [16:0] io_out_0_r_36_im; // @[Reg.scala 19:16]
  reg [16:0] io_out_0_r_37_re; // @[Reg.scala 19:16]
  reg [16:0] io_out_0_r_37_im; // @[Reg.scala 19:16]
  reg [16:0] io_out_0_r_38_re; // @[Reg.scala 19:16]
  reg [16:0] io_out_0_r_38_im; // @[Reg.scala 19:16]
  reg [16:0] io_out_0_r_39_re; // @[Reg.scala 19:16]
  reg [16:0] io_out_0_r_39_im; // @[Reg.scala 19:16]
  reg [16:0] io_out_0_r_40_re; // @[Reg.scala 19:16]
  reg [16:0] io_out_0_r_40_im; // @[Reg.scala 19:16]
  reg [16:0] io_out_0_r_41_re; // @[Reg.scala 19:16]
  reg [16:0] io_out_0_r_41_im; // @[Reg.scala 19:16]
  reg [16:0] io_out_0_r_42_re; // @[Reg.scala 19:16]
  reg [16:0] io_out_0_r_42_im; // @[Reg.scala 19:16]
  reg [16:0] io_out_0_r_43_re; // @[Reg.scala 19:16]
  reg [16:0] io_out_0_r_43_im; // @[Reg.scala 19:16]
  reg [16:0] io_out_0_r_44_re; // @[Reg.scala 19:16]
  reg [16:0] io_out_0_r_44_im; // @[Reg.scala 19:16]
  reg [16:0] io_out_0_r_45_re; // @[Reg.scala 19:16]
  reg [16:0] io_out_0_r_45_im; // @[Reg.scala 19:16]
  reg [16:0] io_out_0_r_46_re; // @[Reg.scala 19:16]
  reg [16:0] io_out_0_r_46_im; // @[Reg.scala 19:16]
  reg [16:0] io_out_0_r_47_re; // @[Reg.scala 19:16]
  reg [16:0] io_out_0_r_47_im; // @[Reg.scala 19:16]
  reg [16:0] io_out_0_r_48_re; // @[Reg.scala 19:16]
  reg [16:0] io_out_0_r_48_im; // @[Reg.scala 19:16]
  reg [16:0] io_out_0_r_49_re; // @[Reg.scala 19:16]
  reg [16:0] io_out_0_r_49_im; // @[Reg.scala 19:16]
  reg [16:0] io_out_0_r_50_re; // @[Reg.scala 19:16]
  reg [16:0] io_out_0_r_50_im; // @[Reg.scala 19:16]
  reg [16:0] io_out_0_r_51_re; // @[Reg.scala 19:16]
  reg [16:0] io_out_0_r_51_im; // @[Reg.scala 19:16]
  reg [16:0] io_out_0_r_52_re; // @[Reg.scala 19:16]
  reg [16:0] io_out_0_r_52_im; // @[Reg.scala 19:16]
  reg [16:0] io_out_0_r_53_re; // @[Reg.scala 19:16]
  reg [16:0] io_out_0_r_53_im; // @[Reg.scala 19:16]
  reg [16:0] io_out_0_r_54_re; // @[Reg.scala 19:16]
  reg [16:0] io_out_0_r_54_im; // @[Reg.scala 19:16]
  reg [16:0] io_out_0_r_55_re; // @[Reg.scala 19:16]
  reg [16:0] io_out_0_r_55_im; // @[Reg.scala 19:16]
  reg [16:0] io_out_0_r_56_re; // @[Reg.scala 19:16]
  reg [16:0] io_out_0_r_56_im; // @[Reg.scala 19:16]
  reg [16:0] io_out_0_r_57_re; // @[Reg.scala 19:16]
  reg [16:0] io_out_0_r_57_im; // @[Reg.scala 19:16]
  reg [16:0] io_out_0_r_58_re; // @[Reg.scala 19:16]
  reg [16:0] io_out_0_r_58_im; // @[Reg.scala 19:16]
  reg [16:0] io_out_0_r_59_re; // @[Reg.scala 19:16]
  reg [16:0] io_out_0_r_59_im; // @[Reg.scala 19:16]
  reg [16:0] io_out_0_r_60_re; // @[Reg.scala 19:16]
  reg [16:0] io_out_0_r_60_im; // @[Reg.scala 19:16]
  reg [16:0] io_out_0_r_61_re; // @[Reg.scala 19:16]
  reg [16:0] io_out_0_r_61_im; // @[Reg.scala 19:16]
  reg [16:0] io_out_0_r_62_re; // @[Reg.scala 19:16]
  reg [16:0] io_out_0_r_62_im; // @[Reg.scala 19:16]
  reg [16:0] io_out_0_r_63_re; // @[Reg.scala 19:16]
  reg [16:0] io_out_0_r_63_im; // @[Reg.scala 19:16]
  assign io_out_0_re = io_out_0_r_63_re; // @[Modules.scala 306:38]
  assign io_out_0_im = io_out_0_r_63_im; // @[Modules.scala 306:38]
  assign io_out_1_re = io_sel ? io_in_0_re : swdata_1_r_63_re; // @[Modules.scala 306:{38,38}]
  assign io_out_1_im = io_sel ? io_in_0_im : swdata_1_r_63_im; // @[Modules.scala 306:{38,38}]
  always @(posedge clock) begin
    swdata_1_r_re <= io_in_1_re; // @[Reg.scala 19:16 20:{18,22}]
    swdata_1_r_im <= io_in_1_im; // @[Reg.scala 19:16 20:{18,22}]
    swdata_1_r_1_re <= swdata_1_r_re; // @[Reg.scala 19:16 20:{18,22}]
    swdata_1_r_1_im <= swdata_1_r_im; // @[Reg.scala 19:16 20:{18,22}]
    swdata_1_r_2_re <= swdata_1_r_1_re; // @[Reg.scala 19:16 20:{18,22}]
    swdata_1_r_2_im <= swdata_1_r_1_im; // @[Reg.scala 19:16 20:{18,22}]
    swdata_1_r_3_re <= swdata_1_r_2_re; // @[Reg.scala 19:16 20:{18,22}]
    swdata_1_r_3_im <= swdata_1_r_2_im; // @[Reg.scala 19:16 20:{18,22}]
    swdata_1_r_4_re <= swdata_1_r_3_re; // @[Reg.scala 19:16 20:{18,22}]
    swdata_1_r_4_im <= swdata_1_r_3_im; // @[Reg.scala 19:16 20:{18,22}]
    swdata_1_r_5_re <= swdata_1_r_4_re; // @[Reg.scala 19:16 20:{18,22}]
    swdata_1_r_5_im <= swdata_1_r_4_im; // @[Reg.scala 19:16 20:{18,22}]
    swdata_1_r_6_re <= swdata_1_r_5_re; // @[Reg.scala 19:16 20:{18,22}]
    swdata_1_r_6_im <= swdata_1_r_5_im; // @[Reg.scala 19:16 20:{18,22}]
    swdata_1_r_7_re <= swdata_1_r_6_re; // @[Reg.scala 19:16 20:{18,22}]
    swdata_1_r_7_im <= swdata_1_r_6_im; // @[Reg.scala 19:16 20:{18,22}]
    swdata_1_r_8_re <= swdata_1_r_7_re; // @[Reg.scala 19:16 20:{18,22}]
    swdata_1_r_8_im <= swdata_1_r_7_im; // @[Reg.scala 19:16 20:{18,22}]
    swdata_1_r_9_re <= swdata_1_r_8_re; // @[Reg.scala 19:16 20:{18,22}]
    swdata_1_r_9_im <= swdata_1_r_8_im; // @[Reg.scala 19:16 20:{18,22}]
    swdata_1_r_10_re <= swdata_1_r_9_re; // @[Reg.scala 19:16 20:{18,22}]
    swdata_1_r_10_im <= swdata_1_r_9_im; // @[Reg.scala 19:16 20:{18,22}]
    swdata_1_r_11_re <= swdata_1_r_10_re; // @[Reg.scala 19:16 20:{18,22}]
    swdata_1_r_11_im <= swdata_1_r_10_im; // @[Reg.scala 19:16 20:{18,22}]
    swdata_1_r_12_re <= swdata_1_r_11_re; // @[Reg.scala 19:16 20:{18,22}]
    swdata_1_r_12_im <= swdata_1_r_11_im; // @[Reg.scala 19:16 20:{18,22}]
    swdata_1_r_13_re <= swdata_1_r_12_re; // @[Reg.scala 19:16 20:{18,22}]
    swdata_1_r_13_im <= swdata_1_r_12_im; // @[Reg.scala 19:16 20:{18,22}]
    swdata_1_r_14_re <= swdata_1_r_13_re; // @[Reg.scala 19:16 20:{18,22}]
    swdata_1_r_14_im <= swdata_1_r_13_im; // @[Reg.scala 19:16 20:{18,22}]
    swdata_1_r_15_re <= swdata_1_r_14_re; // @[Reg.scala 19:16 20:{18,22}]
    swdata_1_r_15_im <= swdata_1_r_14_im; // @[Reg.scala 19:16 20:{18,22}]
    swdata_1_r_16_re <= swdata_1_r_15_re; // @[Reg.scala 19:16 20:{18,22}]
    swdata_1_r_16_im <= swdata_1_r_15_im; // @[Reg.scala 19:16 20:{18,22}]
    swdata_1_r_17_re <= swdata_1_r_16_re; // @[Reg.scala 19:16 20:{18,22}]
    swdata_1_r_17_im <= swdata_1_r_16_im; // @[Reg.scala 19:16 20:{18,22}]
    swdata_1_r_18_re <= swdata_1_r_17_re; // @[Reg.scala 19:16 20:{18,22}]
    swdata_1_r_18_im <= swdata_1_r_17_im; // @[Reg.scala 19:16 20:{18,22}]
    swdata_1_r_19_re <= swdata_1_r_18_re; // @[Reg.scala 19:16 20:{18,22}]
    swdata_1_r_19_im <= swdata_1_r_18_im; // @[Reg.scala 19:16 20:{18,22}]
    swdata_1_r_20_re <= swdata_1_r_19_re; // @[Reg.scala 19:16 20:{18,22}]
    swdata_1_r_20_im <= swdata_1_r_19_im; // @[Reg.scala 19:16 20:{18,22}]
    swdata_1_r_21_re <= swdata_1_r_20_re; // @[Reg.scala 19:16 20:{18,22}]
    swdata_1_r_21_im <= swdata_1_r_20_im; // @[Reg.scala 19:16 20:{18,22}]
    swdata_1_r_22_re <= swdata_1_r_21_re; // @[Reg.scala 19:16 20:{18,22}]
    swdata_1_r_22_im <= swdata_1_r_21_im; // @[Reg.scala 19:16 20:{18,22}]
    swdata_1_r_23_re <= swdata_1_r_22_re; // @[Reg.scala 19:16 20:{18,22}]
    swdata_1_r_23_im <= swdata_1_r_22_im; // @[Reg.scala 19:16 20:{18,22}]
    swdata_1_r_24_re <= swdata_1_r_23_re; // @[Reg.scala 19:16 20:{18,22}]
    swdata_1_r_24_im <= swdata_1_r_23_im; // @[Reg.scala 19:16 20:{18,22}]
    swdata_1_r_25_re <= swdata_1_r_24_re; // @[Reg.scala 19:16 20:{18,22}]
    swdata_1_r_25_im <= swdata_1_r_24_im; // @[Reg.scala 19:16 20:{18,22}]
    swdata_1_r_26_re <= swdata_1_r_25_re; // @[Reg.scala 19:16 20:{18,22}]
    swdata_1_r_26_im <= swdata_1_r_25_im; // @[Reg.scala 19:16 20:{18,22}]
    swdata_1_r_27_re <= swdata_1_r_26_re; // @[Reg.scala 19:16 20:{18,22}]
    swdata_1_r_27_im <= swdata_1_r_26_im; // @[Reg.scala 19:16 20:{18,22}]
    swdata_1_r_28_re <= swdata_1_r_27_re; // @[Reg.scala 19:16 20:{18,22}]
    swdata_1_r_28_im <= swdata_1_r_27_im; // @[Reg.scala 19:16 20:{18,22}]
    swdata_1_r_29_re <= swdata_1_r_28_re; // @[Reg.scala 19:16 20:{18,22}]
    swdata_1_r_29_im <= swdata_1_r_28_im; // @[Reg.scala 19:16 20:{18,22}]
    swdata_1_r_30_re <= swdata_1_r_29_re; // @[Reg.scala 19:16 20:{18,22}]
    swdata_1_r_30_im <= swdata_1_r_29_im; // @[Reg.scala 19:16 20:{18,22}]
    swdata_1_r_31_re <= swdata_1_r_30_re; // @[Reg.scala 19:16 20:{18,22}]
    swdata_1_r_31_im <= swdata_1_r_30_im; // @[Reg.scala 19:16 20:{18,22}]
    swdata_1_r_32_re <= swdata_1_r_31_re; // @[Reg.scala 19:16 20:{18,22}]
    swdata_1_r_32_im <= swdata_1_r_31_im; // @[Reg.scala 19:16 20:{18,22}]
    swdata_1_r_33_re <= swdata_1_r_32_re; // @[Reg.scala 19:16 20:{18,22}]
    swdata_1_r_33_im <= swdata_1_r_32_im; // @[Reg.scala 19:16 20:{18,22}]
    swdata_1_r_34_re <= swdata_1_r_33_re; // @[Reg.scala 19:16 20:{18,22}]
    swdata_1_r_34_im <= swdata_1_r_33_im; // @[Reg.scala 19:16 20:{18,22}]
    swdata_1_r_35_re <= swdata_1_r_34_re; // @[Reg.scala 19:16 20:{18,22}]
    swdata_1_r_35_im <= swdata_1_r_34_im; // @[Reg.scala 19:16 20:{18,22}]
    swdata_1_r_36_re <= swdata_1_r_35_re; // @[Reg.scala 19:16 20:{18,22}]
    swdata_1_r_36_im <= swdata_1_r_35_im; // @[Reg.scala 19:16 20:{18,22}]
    swdata_1_r_37_re <= swdata_1_r_36_re; // @[Reg.scala 19:16 20:{18,22}]
    swdata_1_r_37_im <= swdata_1_r_36_im; // @[Reg.scala 19:16 20:{18,22}]
    swdata_1_r_38_re <= swdata_1_r_37_re; // @[Reg.scala 19:16 20:{18,22}]
    swdata_1_r_38_im <= swdata_1_r_37_im; // @[Reg.scala 19:16 20:{18,22}]
    swdata_1_r_39_re <= swdata_1_r_38_re; // @[Reg.scala 19:16 20:{18,22}]
    swdata_1_r_39_im <= swdata_1_r_38_im; // @[Reg.scala 19:16 20:{18,22}]
    swdata_1_r_40_re <= swdata_1_r_39_re; // @[Reg.scala 19:16 20:{18,22}]
    swdata_1_r_40_im <= swdata_1_r_39_im; // @[Reg.scala 19:16 20:{18,22}]
    swdata_1_r_41_re <= swdata_1_r_40_re; // @[Reg.scala 19:16 20:{18,22}]
    swdata_1_r_41_im <= swdata_1_r_40_im; // @[Reg.scala 19:16 20:{18,22}]
    swdata_1_r_42_re <= swdata_1_r_41_re; // @[Reg.scala 19:16 20:{18,22}]
    swdata_1_r_42_im <= swdata_1_r_41_im; // @[Reg.scala 19:16 20:{18,22}]
    swdata_1_r_43_re <= swdata_1_r_42_re; // @[Reg.scala 19:16 20:{18,22}]
    swdata_1_r_43_im <= swdata_1_r_42_im; // @[Reg.scala 19:16 20:{18,22}]
    swdata_1_r_44_re <= swdata_1_r_43_re; // @[Reg.scala 19:16 20:{18,22}]
    swdata_1_r_44_im <= swdata_1_r_43_im; // @[Reg.scala 19:16 20:{18,22}]
    swdata_1_r_45_re <= swdata_1_r_44_re; // @[Reg.scala 19:16 20:{18,22}]
    swdata_1_r_45_im <= swdata_1_r_44_im; // @[Reg.scala 19:16 20:{18,22}]
    swdata_1_r_46_re <= swdata_1_r_45_re; // @[Reg.scala 19:16 20:{18,22}]
    swdata_1_r_46_im <= swdata_1_r_45_im; // @[Reg.scala 19:16 20:{18,22}]
    swdata_1_r_47_re <= swdata_1_r_46_re; // @[Reg.scala 19:16 20:{18,22}]
    swdata_1_r_47_im <= swdata_1_r_46_im; // @[Reg.scala 19:16 20:{18,22}]
    swdata_1_r_48_re <= swdata_1_r_47_re; // @[Reg.scala 19:16 20:{18,22}]
    swdata_1_r_48_im <= swdata_1_r_47_im; // @[Reg.scala 19:16 20:{18,22}]
    swdata_1_r_49_re <= swdata_1_r_48_re; // @[Reg.scala 19:16 20:{18,22}]
    swdata_1_r_49_im <= swdata_1_r_48_im; // @[Reg.scala 19:16 20:{18,22}]
    swdata_1_r_50_re <= swdata_1_r_49_re; // @[Reg.scala 19:16 20:{18,22}]
    swdata_1_r_50_im <= swdata_1_r_49_im; // @[Reg.scala 19:16 20:{18,22}]
    swdata_1_r_51_re <= swdata_1_r_50_re; // @[Reg.scala 19:16 20:{18,22}]
    swdata_1_r_51_im <= swdata_1_r_50_im; // @[Reg.scala 19:16 20:{18,22}]
    swdata_1_r_52_re <= swdata_1_r_51_re; // @[Reg.scala 19:16 20:{18,22}]
    swdata_1_r_52_im <= swdata_1_r_51_im; // @[Reg.scala 19:16 20:{18,22}]
    swdata_1_r_53_re <= swdata_1_r_52_re; // @[Reg.scala 19:16 20:{18,22}]
    swdata_1_r_53_im <= swdata_1_r_52_im; // @[Reg.scala 19:16 20:{18,22}]
    swdata_1_r_54_re <= swdata_1_r_53_re; // @[Reg.scala 19:16 20:{18,22}]
    swdata_1_r_54_im <= swdata_1_r_53_im; // @[Reg.scala 19:16 20:{18,22}]
    swdata_1_r_55_re <= swdata_1_r_54_re; // @[Reg.scala 19:16 20:{18,22}]
    swdata_1_r_55_im <= swdata_1_r_54_im; // @[Reg.scala 19:16 20:{18,22}]
    swdata_1_r_56_re <= swdata_1_r_55_re; // @[Reg.scala 19:16 20:{18,22}]
    swdata_1_r_56_im <= swdata_1_r_55_im; // @[Reg.scala 19:16 20:{18,22}]
    swdata_1_r_57_re <= swdata_1_r_56_re; // @[Reg.scala 19:16 20:{18,22}]
    swdata_1_r_57_im <= swdata_1_r_56_im; // @[Reg.scala 19:16 20:{18,22}]
    swdata_1_r_58_re <= swdata_1_r_57_re; // @[Reg.scala 19:16 20:{18,22}]
    swdata_1_r_58_im <= swdata_1_r_57_im; // @[Reg.scala 19:16 20:{18,22}]
    swdata_1_r_59_re <= swdata_1_r_58_re; // @[Reg.scala 19:16 20:{18,22}]
    swdata_1_r_59_im <= swdata_1_r_58_im; // @[Reg.scala 19:16 20:{18,22}]
    swdata_1_r_60_re <= swdata_1_r_59_re; // @[Reg.scala 19:16 20:{18,22}]
    swdata_1_r_60_im <= swdata_1_r_59_im; // @[Reg.scala 19:16 20:{18,22}]
    swdata_1_r_61_re <= swdata_1_r_60_re; // @[Reg.scala 19:16 20:{18,22}]
    swdata_1_r_61_im <= swdata_1_r_60_im; // @[Reg.scala 19:16 20:{18,22}]
    swdata_1_r_62_re <= swdata_1_r_61_re; // @[Reg.scala 19:16 20:{18,22}]
    swdata_1_r_62_im <= swdata_1_r_61_im; // @[Reg.scala 19:16 20:{18,22}]
    swdata_1_r_63_re <= swdata_1_r_62_re; // @[Reg.scala 19:16 20:{18,22}]
    swdata_1_r_63_im <= swdata_1_r_62_im; // @[Reg.scala 19:16 20:{18,22}]
    if (io_sel) begin // @[Reg.scala 20:22]
      io_out_0_r_re <= swdata_1_r_63_re; // @[Reg.scala 20:22]
    end else begin
      io_out_0_r_re <= io_in_0_re;
    end
    if (io_sel) begin // @[Reg.scala 20:22]
      io_out_0_r_im <= swdata_1_r_63_im; // @[Reg.scala 20:22]
    end else begin
      io_out_0_r_im <= io_in_0_im;
    end
    io_out_0_r_1_re <= io_out_0_r_re; // @[Reg.scala 19:16 20:{18,22}]
    io_out_0_r_1_im <= io_out_0_r_im; // @[Reg.scala 19:16 20:{18,22}]
    io_out_0_r_2_re <= io_out_0_r_1_re; // @[Reg.scala 19:16 20:{18,22}]
    io_out_0_r_2_im <= io_out_0_r_1_im; // @[Reg.scala 19:16 20:{18,22}]
    io_out_0_r_3_re <= io_out_0_r_2_re; // @[Reg.scala 19:16 20:{18,22}]
    io_out_0_r_3_im <= io_out_0_r_2_im; // @[Reg.scala 19:16 20:{18,22}]
    io_out_0_r_4_re <= io_out_0_r_3_re; // @[Reg.scala 19:16 20:{18,22}]
    io_out_0_r_4_im <= io_out_0_r_3_im; // @[Reg.scala 19:16 20:{18,22}]
    io_out_0_r_5_re <= io_out_0_r_4_re; // @[Reg.scala 19:16 20:{18,22}]
    io_out_0_r_5_im <= io_out_0_r_4_im; // @[Reg.scala 19:16 20:{18,22}]
    io_out_0_r_6_re <= io_out_0_r_5_re; // @[Reg.scala 19:16 20:{18,22}]
    io_out_0_r_6_im <= io_out_0_r_5_im; // @[Reg.scala 19:16 20:{18,22}]
    io_out_0_r_7_re <= io_out_0_r_6_re; // @[Reg.scala 19:16 20:{18,22}]
    io_out_0_r_7_im <= io_out_0_r_6_im; // @[Reg.scala 19:16 20:{18,22}]
    io_out_0_r_8_re <= io_out_0_r_7_re; // @[Reg.scala 19:16 20:{18,22}]
    io_out_0_r_8_im <= io_out_0_r_7_im; // @[Reg.scala 19:16 20:{18,22}]
    io_out_0_r_9_re <= io_out_0_r_8_re; // @[Reg.scala 19:16 20:{18,22}]
    io_out_0_r_9_im <= io_out_0_r_8_im; // @[Reg.scala 19:16 20:{18,22}]
    io_out_0_r_10_re <= io_out_0_r_9_re; // @[Reg.scala 19:16 20:{18,22}]
    io_out_0_r_10_im <= io_out_0_r_9_im; // @[Reg.scala 19:16 20:{18,22}]
    io_out_0_r_11_re <= io_out_0_r_10_re; // @[Reg.scala 19:16 20:{18,22}]
    io_out_0_r_11_im <= io_out_0_r_10_im; // @[Reg.scala 19:16 20:{18,22}]
    io_out_0_r_12_re <= io_out_0_r_11_re; // @[Reg.scala 19:16 20:{18,22}]
    io_out_0_r_12_im <= io_out_0_r_11_im; // @[Reg.scala 19:16 20:{18,22}]
    io_out_0_r_13_re <= io_out_0_r_12_re; // @[Reg.scala 19:16 20:{18,22}]
    io_out_0_r_13_im <= io_out_0_r_12_im; // @[Reg.scala 19:16 20:{18,22}]
    io_out_0_r_14_re <= io_out_0_r_13_re; // @[Reg.scala 19:16 20:{18,22}]
    io_out_0_r_14_im <= io_out_0_r_13_im; // @[Reg.scala 19:16 20:{18,22}]
    io_out_0_r_15_re <= io_out_0_r_14_re; // @[Reg.scala 19:16 20:{18,22}]
    io_out_0_r_15_im <= io_out_0_r_14_im; // @[Reg.scala 19:16 20:{18,22}]
    io_out_0_r_16_re <= io_out_0_r_15_re; // @[Reg.scala 19:16 20:{18,22}]
    io_out_0_r_16_im <= io_out_0_r_15_im; // @[Reg.scala 19:16 20:{18,22}]
    io_out_0_r_17_re <= io_out_0_r_16_re; // @[Reg.scala 19:16 20:{18,22}]
    io_out_0_r_17_im <= io_out_0_r_16_im; // @[Reg.scala 19:16 20:{18,22}]
    io_out_0_r_18_re <= io_out_0_r_17_re; // @[Reg.scala 19:16 20:{18,22}]
    io_out_0_r_18_im <= io_out_0_r_17_im; // @[Reg.scala 19:16 20:{18,22}]
    io_out_0_r_19_re <= io_out_0_r_18_re; // @[Reg.scala 19:16 20:{18,22}]
    io_out_0_r_19_im <= io_out_0_r_18_im; // @[Reg.scala 19:16 20:{18,22}]
    io_out_0_r_20_re <= io_out_0_r_19_re; // @[Reg.scala 19:16 20:{18,22}]
    io_out_0_r_20_im <= io_out_0_r_19_im; // @[Reg.scala 19:16 20:{18,22}]
    io_out_0_r_21_re <= io_out_0_r_20_re; // @[Reg.scala 19:16 20:{18,22}]
    io_out_0_r_21_im <= io_out_0_r_20_im; // @[Reg.scala 19:16 20:{18,22}]
    io_out_0_r_22_re <= io_out_0_r_21_re; // @[Reg.scala 19:16 20:{18,22}]
    io_out_0_r_22_im <= io_out_0_r_21_im; // @[Reg.scala 19:16 20:{18,22}]
    io_out_0_r_23_re <= io_out_0_r_22_re; // @[Reg.scala 19:16 20:{18,22}]
    io_out_0_r_23_im <= io_out_0_r_22_im; // @[Reg.scala 19:16 20:{18,22}]
    io_out_0_r_24_re <= io_out_0_r_23_re; // @[Reg.scala 19:16 20:{18,22}]
    io_out_0_r_24_im <= io_out_0_r_23_im; // @[Reg.scala 19:16 20:{18,22}]
    io_out_0_r_25_re <= io_out_0_r_24_re; // @[Reg.scala 19:16 20:{18,22}]
    io_out_0_r_25_im <= io_out_0_r_24_im; // @[Reg.scala 19:16 20:{18,22}]
    io_out_0_r_26_re <= io_out_0_r_25_re; // @[Reg.scala 19:16 20:{18,22}]
    io_out_0_r_26_im <= io_out_0_r_25_im; // @[Reg.scala 19:16 20:{18,22}]
    io_out_0_r_27_re <= io_out_0_r_26_re; // @[Reg.scala 19:16 20:{18,22}]
    io_out_0_r_27_im <= io_out_0_r_26_im; // @[Reg.scala 19:16 20:{18,22}]
    io_out_0_r_28_re <= io_out_0_r_27_re; // @[Reg.scala 19:16 20:{18,22}]
    io_out_0_r_28_im <= io_out_0_r_27_im; // @[Reg.scala 19:16 20:{18,22}]
    io_out_0_r_29_re <= io_out_0_r_28_re; // @[Reg.scala 19:16 20:{18,22}]
    io_out_0_r_29_im <= io_out_0_r_28_im; // @[Reg.scala 19:16 20:{18,22}]
    io_out_0_r_30_re <= io_out_0_r_29_re; // @[Reg.scala 19:16 20:{18,22}]
    io_out_0_r_30_im <= io_out_0_r_29_im; // @[Reg.scala 19:16 20:{18,22}]
    io_out_0_r_31_re <= io_out_0_r_30_re; // @[Reg.scala 19:16 20:{18,22}]
    io_out_0_r_31_im <= io_out_0_r_30_im; // @[Reg.scala 19:16 20:{18,22}]
    io_out_0_r_32_re <= io_out_0_r_31_re; // @[Reg.scala 19:16 20:{18,22}]
    io_out_0_r_32_im <= io_out_0_r_31_im; // @[Reg.scala 19:16 20:{18,22}]
    io_out_0_r_33_re <= io_out_0_r_32_re; // @[Reg.scala 19:16 20:{18,22}]
    io_out_0_r_33_im <= io_out_0_r_32_im; // @[Reg.scala 19:16 20:{18,22}]
    io_out_0_r_34_re <= io_out_0_r_33_re; // @[Reg.scala 19:16 20:{18,22}]
    io_out_0_r_34_im <= io_out_0_r_33_im; // @[Reg.scala 19:16 20:{18,22}]
    io_out_0_r_35_re <= io_out_0_r_34_re; // @[Reg.scala 19:16 20:{18,22}]
    io_out_0_r_35_im <= io_out_0_r_34_im; // @[Reg.scala 19:16 20:{18,22}]
    io_out_0_r_36_re <= io_out_0_r_35_re; // @[Reg.scala 19:16 20:{18,22}]
    io_out_0_r_36_im <= io_out_0_r_35_im; // @[Reg.scala 19:16 20:{18,22}]
    io_out_0_r_37_re <= io_out_0_r_36_re; // @[Reg.scala 19:16 20:{18,22}]
    io_out_0_r_37_im <= io_out_0_r_36_im; // @[Reg.scala 19:16 20:{18,22}]
    io_out_0_r_38_re <= io_out_0_r_37_re; // @[Reg.scala 19:16 20:{18,22}]
    io_out_0_r_38_im <= io_out_0_r_37_im; // @[Reg.scala 19:16 20:{18,22}]
    io_out_0_r_39_re <= io_out_0_r_38_re; // @[Reg.scala 19:16 20:{18,22}]
    io_out_0_r_39_im <= io_out_0_r_38_im; // @[Reg.scala 19:16 20:{18,22}]
    io_out_0_r_40_re <= io_out_0_r_39_re; // @[Reg.scala 19:16 20:{18,22}]
    io_out_0_r_40_im <= io_out_0_r_39_im; // @[Reg.scala 19:16 20:{18,22}]
    io_out_0_r_41_re <= io_out_0_r_40_re; // @[Reg.scala 19:16 20:{18,22}]
    io_out_0_r_41_im <= io_out_0_r_40_im; // @[Reg.scala 19:16 20:{18,22}]
    io_out_0_r_42_re <= io_out_0_r_41_re; // @[Reg.scala 19:16 20:{18,22}]
    io_out_0_r_42_im <= io_out_0_r_41_im; // @[Reg.scala 19:16 20:{18,22}]
    io_out_0_r_43_re <= io_out_0_r_42_re; // @[Reg.scala 19:16 20:{18,22}]
    io_out_0_r_43_im <= io_out_0_r_42_im; // @[Reg.scala 19:16 20:{18,22}]
    io_out_0_r_44_re <= io_out_0_r_43_re; // @[Reg.scala 19:16 20:{18,22}]
    io_out_0_r_44_im <= io_out_0_r_43_im; // @[Reg.scala 19:16 20:{18,22}]
    io_out_0_r_45_re <= io_out_0_r_44_re; // @[Reg.scala 19:16 20:{18,22}]
    io_out_0_r_45_im <= io_out_0_r_44_im; // @[Reg.scala 19:16 20:{18,22}]
    io_out_0_r_46_re <= io_out_0_r_45_re; // @[Reg.scala 19:16 20:{18,22}]
    io_out_0_r_46_im <= io_out_0_r_45_im; // @[Reg.scala 19:16 20:{18,22}]
    io_out_0_r_47_re <= io_out_0_r_46_re; // @[Reg.scala 19:16 20:{18,22}]
    io_out_0_r_47_im <= io_out_0_r_46_im; // @[Reg.scala 19:16 20:{18,22}]
    io_out_0_r_48_re <= io_out_0_r_47_re; // @[Reg.scala 19:16 20:{18,22}]
    io_out_0_r_48_im <= io_out_0_r_47_im; // @[Reg.scala 19:16 20:{18,22}]
    io_out_0_r_49_re <= io_out_0_r_48_re; // @[Reg.scala 19:16 20:{18,22}]
    io_out_0_r_49_im <= io_out_0_r_48_im; // @[Reg.scala 19:16 20:{18,22}]
    io_out_0_r_50_re <= io_out_0_r_49_re; // @[Reg.scala 19:16 20:{18,22}]
    io_out_0_r_50_im <= io_out_0_r_49_im; // @[Reg.scala 19:16 20:{18,22}]
    io_out_0_r_51_re <= io_out_0_r_50_re; // @[Reg.scala 19:16 20:{18,22}]
    io_out_0_r_51_im <= io_out_0_r_50_im; // @[Reg.scala 19:16 20:{18,22}]
    io_out_0_r_52_re <= io_out_0_r_51_re; // @[Reg.scala 19:16 20:{18,22}]
    io_out_0_r_52_im <= io_out_0_r_51_im; // @[Reg.scala 19:16 20:{18,22}]
    io_out_0_r_53_re <= io_out_0_r_52_re; // @[Reg.scala 19:16 20:{18,22}]
    io_out_0_r_53_im <= io_out_0_r_52_im; // @[Reg.scala 19:16 20:{18,22}]
    io_out_0_r_54_re <= io_out_0_r_53_re; // @[Reg.scala 19:16 20:{18,22}]
    io_out_0_r_54_im <= io_out_0_r_53_im; // @[Reg.scala 19:16 20:{18,22}]
    io_out_0_r_55_re <= io_out_0_r_54_re; // @[Reg.scala 19:16 20:{18,22}]
    io_out_0_r_55_im <= io_out_0_r_54_im; // @[Reg.scala 19:16 20:{18,22}]
    io_out_0_r_56_re <= io_out_0_r_55_re; // @[Reg.scala 19:16 20:{18,22}]
    io_out_0_r_56_im <= io_out_0_r_55_im; // @[Reg.scala 19:16 20:{18,22}]
    io_out_0_r_57_re <= io_out_0_r_56_re; // @[Reg.scala 19:16 20:{18,22}]
    io_out_0_r_57_im <= io_out_0_r_56_im; // @[Reg.scala 19:16 20:{18,22}]
    io_out_0_r_58_re <= io_out_0_r_57_re; // @[Reg.scala 19:16 20:{18,22}]
    io_out_0_r_58_im <= io_out_0_r_57_im; // @[Reg.scala 19:16 20:{18,22}]
    io_out_0_r_59_re <= io_out_0_r_58_re; // @[Reg.scala 19:16 20:{18,22}]
    io_out_0_r_59_im <= io_out_0_r_58_im; // @[Reg.scala 19:16 20:{18,22}]
    io_out_0_r_60_re <= io_out_0_r_59_re; // @[Reg.scala 19:16 20:{18,22}]
    io_out_0_r_60_im <= io_out_0_r_59_im; // @[Reg.scala 19:16 20:{18,22}]
    io_out_0_r_61_re <= io_out_0_r_60_re; // @[Reg.scala 19:16 20:{18,22}]
    io_out_0_r_61_im <= io_out_0_r_60_im; // @[Reg.scala 19:16 20:{18,22}]
    io_out_0_r_62_re <= io_out_0_r_61_re; // @[Reg.scala 19:16 20:{18,22}]
    io_out_0_r_62_im <= io_out_0_r_61_im; // @[Reg.scala 19:16 20:{18,22}]
    io_out_0_r_63_re <= io_out_0_r_62_re; // @[Reg.scala 19:16 20:{18,22}]
    io_out_0_r_63_im <= io_out_0_r_62_im; // @[Reg.scala 19:16 20:{18,22}]
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  swdata_1_r_re = _RAND_0[16:0];
  _RAND_1 = {1{`RANDOM}};
  swdata_1_r_im = _RAND_1[16:0];
  _RAND_2 = {1{`RANDOM}};
  swdata_1_r_1_re = _RAND_2[16:0];
  _RAND_3 = {1{`RANDOM}};
  swdata_1_r_1_im = _RAND_3[16:0];
  _RAND_4 = {1{`RANDOM}};
  swdata_1_r_2_re = _RAND_4[16:0];
  _RAND_5 = {1{`RANDOM}};
  swdata_1_r_2_im = _RAND_5[16:0];
  _RAND_6 = {1{`RANDOM}};
  swdata_1_r_3_re = _RAND_6[16:0];
  _RAND_7 = {1{`RANDOM}};
  swdata_1_r_3_im = _RAND_7[16:0];
  _RAND_8 = {1{`RANDOM}};
  swdata_1_r_4_re = _RAND_8[16:0];
  _RAND_9 = {1{`RANDOM}};
  swdata_1_r_4_im = _RAND_9[16:0];
  _RAND_10 = {1{`RANDOM}};
  swdata_1_r_5_re = _RAND_10[16:0];
  _RAND_11 = {1{`RANDOM}};
  swdata_1_r_5_im = _RAND_11[16:0];
  _RAND_12 = {1{`RANDOM}};
  swdata_1_r_6_re = _RAND_12[16:0];
  _RAND_13 = {1{`RANDOM}};
  swdata_1_r_6_im = _RAND_13[16:0];
  _RAND_14 = {1{`RANDOM}};
  swdata_1_r_7_re = _RAND_14[16:0];
  _RAND_15 = {1{`RANDOM}};
  swdata_1_r_7_im = _RAND_15[16:0];
  _RAND_16 = {1{`RANDOM}};
  swdata_1_r_8_re = _RAND_16[16:0];
  _RAND_17 = {1{`RANDOM}};
  swdata_1_r_8_im = _RAND_17[16:0];
  _RAND_18 = {1{`RANDOM}};
  swdata_1_r_9_re = _RAND_18[16:0];
  _RAND_19 = {1{`RANDOM}};
  swdata_1_r_9_im = _RAND_19[16:0];
  _RAND_20 = {1{`RANDOM}};
  swdata_1_r_10_re = _RAND_20[16:0];
  _RAND_21 = {1{`RANDOM}};
  swdata_1_r_10_im = _RAND_21[16:0];
  _RAND_22 = {1{`RANDOM}};
  swdata_1_r_11_re = _RAND_22[16:0];
  _RAND_23 = {1{`RANDOM}};
  swdata_1_r_11_im = _RAND_23[16:0];
  _RAND_24 = {1{`RANDOM}};
  swdata_1_r_12_re = _RAND_24[16:0];
  _RAND_25 = {1{`RANDOM}};
  swdata_1_r_12_im = _RAND_25[16:0];
  _RAND_26 = {1{`RANDOM}};
  swdata_1_r_13_re = _RAND_26[16:0];
  _RAND_27 = {1{`RANDOM}};
  swdata_1_r_13_im = _RAND_27[16:0];
  _RAND_28 = {1{`RANDOM}};
  swdata_1_r_14_re = _RAND_28[16:0];
  _RAND_29 = {1{`RANDOM}};
  swdata_1_r_14_im = _RAND_29[16:0];
  _RAND_30 = {1{`RANDOM}};
  swdata_1_r_15_re = _RAND_30[16:0];
  _RAND_31 = {1{`RANDOM}};
  swdata_1_r_15_im = _RAND_31[16:0];
  _RAND_32 = {1{`RANDOM}};
  swdata_1_r_16_re = _RAND_32[16:0];
  _RAND_33 = {1{`RANDOM}};
  swdata_1_r_16_im = _RAND_33[16:0];
  _RAND_34 = {1{`RANDOM}};
  swdata_1_r_17_re = _RAND_34[16:0];
  _RAND_35 = {1{`RANDOM}};
  swdata_1_r_17_im = _RAND_35[16:0];
  _RAND_36 = {1{`RANDOM}};
  swdata_1_r_18_re = _RAND_36[16:0];
  _RAND_37 = {1{`RANDOM}};
  swdata_1_r_18_im = _RAND_37[16:0];
  _RAND_38 = {1{`RANDOM}};
  swdata_1_r_19_re = _RAND_38[16:0];
  _RAND_39 = {1{`RANDOM}};
  swdata_1_r_19_im = _RAND_39[16:0];
  _RAND_40 = {1{`RANDOM}};
  swdata_1_r_20_re = _RAND_40[16:0];
  _RAND_41 = {1{`RANDOM}};
  swdata_1_r_20_im = _RAND_41[16:0];
  _RAND_42 = {1{`RANDOM}};
  swdata_1_r_21_re = _RAND_42[16:0];
  _RAND_43 = {1{`RANDOM}};
  swdata_1_r_21_im = _RAND_43[16:0];
  _RAND_44 = {1{`RANDOM}};
  swdata_1_r_22_re = _RAND_44[16:0];
  _RAND_45 = {1{`RANDOM}};
  swdata_1_r_22_im = _RAND_45[16:0];
  _RAND_46 = {1{`RANDOM}};
  swdata_1_r_23_re = _RAND_46[16:0];
  _RAND_47 = {1{`RANDOM}};
  swdata_1_r_23_im = _RAND_47[16:0];
  _RAND_48 = {1{`RANDOM}};
  swdata_1_r_24_re = _RAND_48[16:0];
  _RAND_49 = {1{`RANDOM}};
  swdata_1_r_24_im = _RAND_49[16:0];
  _RAND_50 = {1{`RANDOM}};
  swdata_1_r_25_re = _RAND_50[16:0];
  _RAND_51 = {1{`RANDOM}};
  swdata_1_r_25_im = _RAND_51[16:0];
  _RAND_52 = {1{`RANDOM}};
  swdata_1_r_26_re = _RAND_52[16:0];
  _RAND_53 = {1{`RANDOM}};
  swdata_1_r_26_im = _RAND_53[16:0];
  _RAND_54 = {1{`RANDOM}};
  swdata_1_r_27_re = _RAND_54[16:0];
  _RAND_55 = {1{`RANDOM}};
  swdata_1_r_27_im = _RAND_55[16:0];
  _RAND_56 = {1{`RANDOM}};
  swdata_1_r_28_re = _RAND_56[16:0];
  _RAND_57 = {1{`RANDOM}};
  swdata_1_r_28_im = _RAND_57[16:0];
  _RAND_58 = {1{`RANDOM}};
  swdata_1_r_29_re = _RAND_58[16:0];
  _RAND_59 = {1{`RANDOM}};
  swdata_1_r_29_im = _RAND_59[16:0];
  _RAND_60 = {1{`RANDOM}};
  swdata_1_r_30_re = _RAND_60[16:0];
  _RAND_61 = {1{`RANDOM}};
  swdata_1_r_30_im = _RAND_61[16:0];
  _RAND_62 = {1{`RANDOM}};
  swdata_1_r_31_re = _RAND_62[16:0];
  _RAND_63 = {1{`RANDOM}};
  swdata_1_r_31_im = _RAND_63[16:0];
  _RAND_64 = {1{`RANDOM}};
  swdata_1_r_32_re = _RAND_64[16:0];
  _RAND_65 = {1{`RANDOM}};
  swdata_1_r_32_im = _RAND_65[16:0];
  _RAND_66 = {1{`RANDOM}};
  swdata_1_r_33_re = _RAND_66[16:0];
  _RAND_67 = {1{`RANDOM}};
  swdata_1_r_33_im = _RAND_67[16:0];
  _RAND_68 = {1{`RANDOM}};
  swdata_1_r_34_re = _RAND_68[16:0];
  _RAND_69 = {1{`RANDOM}};
  swdata_1_r_34_im = _RAND_69[16:0];
  _RAND_70 = {1{`RANDOM}};
  swdata_1_r_35_re = _RAND_70[16:0];
  _RAND_71 = {1{`RANDOM}};
  swdata_1_r_35_im = _RAND_71[16:0];
  _RAND_72 = {1{`RANDOM}};
  swdata_1_r_36_re = _RAND_72[16:0];
  _RAND_73 = {1{`RANDOM}};
  swdata_1_r_36_im = _RAND_73[16:0];
  _RAND_74 = {1{`RANDOM}};
  swdata_1_r_37_re = _RAND_74[16:0];
  _RAND_75 = {1{`RANDOM}};
  swdata_1_r_37_im = _RAND_75[16:0];
  _RAND_76 = {1{`RANDOM}};
  swdata_1_r_38_re = _RAND_76[16:0];
  _RAND_77 = {1{`RANDOM}};
  swdata_1_r_38_im = _RAND_77[16:0];
  _RAND_78 = {1{`RANDOM}};
  swdata_1_r_39_re = _RAND_78[16:0];
  _RAND_79 = {1{`RANDOM}};
  swdata_1_r_39_im = _RAND_79[16:0];
  _RAND_80 = {1{`RANDOM}};
  swdata_1_r_40_re = _RAND_80[16:0];
  _RAND_81 = {1{`RANDOM}};
  swdata_1_r_40_im = _RAND_81[16:0];
  _RAND_82 = {1{`RANDOM}};
  swdata_1_r_41_re = _RAND_82[16:0];
  _RAND_83 = {1{`RANDOM}};
  swdata_1_r_41_im = _RAND_83[16:0];
  _RAND_84 = {1{`RANDOM}};
  swdata_1_r_42_re = _RAND_84[16:0];
  _RAND_85 = {1{`RANDOM}};
  swdata_1_r_42_im = _RAND_85[16:0];
  _RAND_86 = {1{`RANDOM}};
  swdata_1_r_43_re = _RAND_86[16:0];
  _RAND_87 = {1{`RANDOM}};
  swdata_1_r_43_im = _RAND_87[16:0];
  _RAND_88 = {1{`RANDOM}};
  swdata_1_r_44_re = _RAND_88[16:0];
  _RAND_89 = {1{`RANDOM}};
  swdata_1_r_44_im = _RAND_89[16:0];
  _RAND_90 = {1{`RANDOM}};
  swdata_1_r_45_re = _RAND_90[16:0];
  _RAND_91 = {1{`RANDOM}};
  swdata_1_r_45_im = _RAND_91[16:0];
  _RAND_92 = {1{`RANDOM}};
  swdata_1_r_46_re = _RAND_92[16:0];
  _RAND_93 = {1{`RANDOM}};
  swdata_1_r_46_im = _RAND_93[16:0];
  _RAND_94 = {1{`RANDOM}};
  swdata_1_r_47_re = _RAND_94[16:0];
  _RAND_95 = {1{`RANDOM}};
  swdata_1_r_47_im = _RAND_95[16:0];
  _RAND_96 = {1{`RANDOM}};
  swdata_1_r_48_re = _RAND_96[16:0];
  _RAND_97 = {1{`RANDOM}};
  swdata_1_r_48_im = _RAND_97[16:0];
  _RAND_98 = {1{`RANDOM}};
  swdata_1_r_49_re = _RAND_98[16:0];
  _RAND_99 = {1{`RANDOM}};
  swdata_1_r_49_im = _RAND_99[16:0];
  _RAND_100 = {1{`RANDOM}};
  swdata_1_r_50_re = _RAND_100[16:0];
  _RAND_101 = {1{`RANDOM}};
  swdata_1_r_50_im = _RAND_101[16:0];
  _RAND_102 = {1{`RANDOM}};
  swdata_1_r_51_re = _RAND_102[16:0];
  _RAND_103 = {1{`RANDOM}};
  swdata_1_r_51_im = _RAND_103[16:0];
  _RAND_104 = {1{`RANDOM}};
  swdata_1_r_52_re = _RAND_104[16:0];
  _RAND_105 = {1{`RANDOM}};
  swdata_1_r_52_im = _RAND_105[16:0];
  _RAND_106 = {1{`RANDOM}};
  swdata_1_r_53_re = _RAND_106[16:0];
  _RAND_107 = {1{`RANDOM}};
  swdata_1_r_53_im = _RAND_107[16:0];
  _RAND_108 = {1{`RANDOM}};
  swdata_1_r_54_re = _RAND_108[16:0];
  _RAND_109 = {1{`RANDOM}};
  swdata_1_r_54_im = _RAND_109[16:0];
  _RAND_110 = {1{`RANDOM}};
  swdata_1_r_55_re = _RAND_110[16:0];
  _RAND_111 = {1{`RANDOM}};
  swdata_1_r_55_im = _RAND_111[16:0];
  _RAND_112 = {1{`RANDOM}};
  swdata_1_r_56_re = _RAND_112[16:0];
  _RAND_113 = {1{`RANDOM}};
  swdata_1_r_56_im = _RAND_113[16:0];
  _RAND_114 = {1{`RANDOM}};
  swdata_1_r_57_re = _RAND_114[16:0];
  _RAND_115 = {1{`RANDOM}};
  swdata_1_r_57_im = _RAND_115[16:0];
  _RAND_116 = {1{`RANDOM}};
  swdata_1_r_58_re = _RAND_116[16:0];
  _RAND_117 = {1{`RANDOM}};
  swdata_1_r_58_im = _RAND_117[16:0];
  _RAND_118 = {1{`RANDOM}};
  swdata_1_r_59_re = _RAND_118[16:0];
  _RAND_119 = {1{`RANDOM}};
  swdata_1_r_59_im = _RAND_119[16:0];
  _RAND_120 = {1{`RANDOM}};
  swdata_1_r_60_re = _RAND_120[16:0];
  _RAND_121 = {1{`RANDOM}};
  swdata_1_r_60_im = _RAND_121[16:0];
  _RAND_122 = {1{`RANDOM}};
  swdata_1_r_61_re = _RAND_122[16:0];
  _RAND_123 = {1{`RANDOM}};
  swdata_1_r_61_im = _RAND_123[16:0];
  _RAND_124 = {1{`RANDOM}};
  swdata_1_r_62_re = _RAND_124[16:0];
  _RAND_125 = {1{`RANDOM}};
  swdata_1_r_62_im = _RAND_125[16:0];
  _RAND_126 = {1{`RANDOM}};
  swdata_1_r_63_re = _RAND_126[16:0];
  _RAND_127 = {1{`RANDOM}};
  swdata_1_r_63_im = _RAND_127[16:0];
  _RAND_128 = {1{`RANDOM}};
  io_out_0_r_re = _RAND_128[16:0];
  _RAND_129 = {1{`RANDOM}};
  io_out_0_r_im = _RAND_129[16:0];
  _RAND_130 = {1{`RANDOM}};
  io_out_0_r_1_re = _RAND_130[16:0];
  _RAND_131 = {1{`RANDOM}};
  io_out_0_r_1_im = _RAND_131[16:0];
  _RAND_132 = {1{`RANDOM}};
  io_out_0_r_2_re = _RAND_132[16:0];
  _RAND_133 = {1{`RANDOM}};
  io_out_0_r_2_im = _RAND_133[16:0];
  _RAND_134 = {1{`RANDOM}};
  io_out_0_r_3_re = _RAND_134[16:0];
  _RAND_135 = {1{`RANDOM}};
  io_out_0_r_3_im = _RAND_135[16:0];
  _RAND_136 = {1{`RANDOM}};
  io_out_0_r_4_re = _RAND_136[16:0];
  _RAND_137 = {1{`RANDOM}};
  io_out_0_r_4_im = _RAND_137[16:0];
  _RAND_138 = {1{`RANDOM}};
  io_out_0_r_5_re = _RAND_138[16:0];
  _RAND_139 = {1{`RANDOM}};
  io_out_0_r_5_im = _RAND_139[16:0];
  _RAND_140 = {1{`RANDOM}};
  io_out_0_r_6_re = _RAND_140[16:0];
  _RAND_141 = {1{`RANDOM}};
  io_out_0_r_6_im = _RAND_141[16:0];
  _RAND_142 = {1{`RANDOM}};
  io_out_0_r_7_re = _RAND_142[16:0];
  _RAND_143 = {1{`RANDOM}};
  io_out_0_r_7_im = _RAND_143[16:0];
  _RAND_144 = {1{`RANDOM}};
  io_out_0_r_8_re = _RAND_144[16:0];
  _RAND_145 = {1{`RANDOM}};
  io_out_0_r_8_im = _RAND_145[16:0];
  _RAND_146 = {1{`RANDOM}};
  io_out_0_r_9_re = _RAND_146[16:0];
  _RAND_147 = {1{`RANDOM}};
  io_out_0_r_9_im = _RAND_147[16:0];
  _RAND_148 = {1{`RANDOM}};
  io_out_0_r_10_re = _RAND_148[16:0];
  _RAND_149 = {1{`RANDOM}};
  io_out_0_r_10_im = _RAND_149[16:0];
  _RAND_150 = {1{`RANDOM}};
  io_out_0_r_11_re = _RAND_150[16:0];
  _RAND_151 = {1{`RANDOM}};
  io_out_0_r_11_im = _RAND_151[16:0];
  _RAND_152 = {1{`RANDOM}};
  io_out_0_r_12_re = _RAND_152[16:0];
  _RAND_153 = {1{`RANDOM}};
  io_out_0_r_12_im = _RAND_153[16:0];
  _RAND_154 = {1{`RANDOM}};
  io_out_0_r_13_re = _RAND_154[16:0];
  _RAND_155 = {1{`RANDOM}};
  io_out_0_r_13_im = _RAND_155[16:0];
  _RAND_156 = {1{`RANDOM}};
  io_out_0_r_14_re = _RAND_156[16:0];
  _RAND_157 = {1{`RANDOM}};
  io_out_0_r_14_im = _RAND_157[16:0];
  _RAND_158 = {1{`RANDOM}};
  io_out_0_r_15_re = _RAND_158[16:0];
  _RAND_159 = {1{`RANDOM}};
  io_out_0_r_15_im = _RAND_159[16:0];
  _RAND_160 = {1{`RANDOM}};
  io_out_0_r_16_re = _RAND_160[16:0];
  _RAND_161 = {1{`RANDOM}};
  io_out_0_r_16_im = _RAND_161[16:0];
  _RAND_162 = {1{`RANDOM}};
  io_out_0_r_17_re = _RAND_162[16:0];
  _RAND_163 = {1{`RANDOM}};
  io_out_0_r_17_im = _RAND_163[16:0];
  _RAND_164 = {1{`RANDOM}};
  io_out_0_r_18_re = _RAND_164[16:0];
  _RAND_165 = {1{`RANDOM}};
  io_out_0_r_18_im = _RAND_165[16:0];
  _RAND_166 = {1{`RANDOM}};
  io_out_0_r_19_re = _RAND_166[16:0];
  _RAND_167 = {1{`RANDOM}};
  io_out_0_r_19_im = _RAND_167[16:0];
  _RAND_168 = {1{`RANDOM}};
  io_out_0_r_20_re = _RAND_168[16:0];
  _RAND_169 = {1{`RANDOM}};
  io_out_0_r_20_im = _RAND_169[16:0];
  _RAND_170 = {1{`RANDOM}};
  io_out_0_r_21_re = _RAND_170[16:0];
  _RAND_171 = {1{`RANDOM}};
  io_out_0_r_21_im = _RAND_171[16:0];
  _RAND_172 = {1{`RANDOM}};
  io_out_0_r_22_re = _RAND_172[16:0];
  _RAND_173 = {1{`RANDOM}};
  io_out_0_r_22_im = _RAND_173[16:0];
  _RAND_174 = {1{`RANDOM}};
  io_out_0_r_23_re = _RAND_174[16:0];
  _RAND_175 = {1{`RANDOM}};
  io_out_0_r_23_im = _RAND_175[16:0];
  _RAND_176 = {1{`RANDOM}};
  io_out_0_r_24_re = _RAND_176[16:0];
  _RAND_177 = {1{`RANDOM}};
  io_out_0_r_24_im = _RAND_177[16:0];
  _RAND_178 = {1{`RANDOM}};
  io_out_0_r_25_re = _RAND_178[16:0];
  _RAND_179 = {1{`RANDOM}};
  io_out_0_r_25_im = _RAND_179[16:0];
  _RAND_180 = {1{`RANDOM}};
  io_out_0_r_26_re = _RAND_180[16:0];
  _RAND_181 = {1{`RANDOM}};
  io_out_0_r_26_im = _RAND_181[16:0];
  _RAND_182 = {1{`RANDOM}};
  io_out_0_r_27_re = _RAND_182[16:0];
  _RAND_183 = {1{`RANDOM}};
  io_out_0_r_27_im = _RAND_183[16:0];
  _RAND_184 = {1{`RANDOM}};
  io_out_0_r_28_re = _RAND_184[16:0];
  _RAND_185 = {1{`RANDOM}};
  io_out_0_r_28_im = _RAND_185[16:0];
  _RAND_186 = {1{`RANDOM}};
  io_out_0_r_29_re = _RAND_186[16:0];
  _RAND_187 = {1{`RANDOM}};
  io_out_0_r_29_im = _RAND_187[16:0];
  _RAND_188 = {1{`RANDOM}};
  io_out_0_r_30_re = _RAND_188[16:0];
  _RAND_189 = {1{`RANDOM}};
  io_out_0_r_30_im = _RAND_189[16:0];
  _RAND_190 = {1{`RANDOM}};
  io_out_0_r_31_re = _RAND_190[16:0];
  _RAND_191 = {1{`RANDOM}};
  io_out_0_r_31_im = _RAND_191[16:0];
  _RAND_192 = {1{`RANDOM}};
  io_out_0_r_32_re = _RAND_192[16:0];
  _RAND_193 = {1{`RANDOM}};
  io_out_0_r_32_im = _RAND_193[16:0];
  _RAND_194 = {1{`RANDOM}};
  io_out_0_r_33_re = _RAND_194[16:0];
  _RAND_195 = {1{`RANDOM}};
  io_out_0_r_33_im = _RAND_195[16:0];
  _RAND_196 = {1{`RANDOM}};
  io_out_0_r_34_re = _RAND_196[16:0];
  _RAND_197 = {1{`RANDOM}};
  io_out_0_r_34_im = _RAND_197[16:0];
  _RAND_198 = {1{`RANDOM}};
  io_out_0_r_35_re = _RAND_198[16:0];
  _RAND_199 = {1{`RANDOM}};
  io_out_0_r_35_im = _RAND_199[16:0];
  _RAND_200 = {1{`RANDOM}};
  io_out_0_r_36_re = _RAND_200[16:0];
  _RAND_201 = {1{`RANDOM}};
  io_out_0_r_36_im = _RAND_201[16:0];
  _RAND_202 = {1{`RANDOM}};
  io_out_0_r_37_re = _RAND_202[16:0];
  _RAND_203 = {1{`RANDOM}};
  io_out_0_r_37_im = _RAND_203[16:0];
  _RAND_204 = {1{`RANDOM}};
  io_out_0_r_38_re = _RAND_204[16:0];
  _RAND_205 = {1{`RANDOM}};
  io_out_0_r_38_im = _RAND_205[16:0];
  _RAND_206 = {1{`RANDOM}};
  io_out_0_r_39_re = _RAND_206[16:0];
  _RAND_207 = {1{`RANDOM}};
  io_out_0_r_39_im = _RAND_207[16:0];
  _RAND_208 = {1{`RANDOM}};
  io_out_0_r_40_re = _RAND_208[16:0];
  _RAND_209 = {1{`RANDOM}};
  io_out_0_r_40_im = _RAND_209[16:0];
  _RAND_210 = {1{`RANDOM}};
  io_out_0_r_41_re = _RAND_210[16:0];
  _RAND_211 = {1{`RANDOM}};
  io_out_0_r_41_im = _RAND_211[16:0];
  _RAND_212 = {1{`RANDOM}};
  io_out_0_r_42_re = _RAND_212[16:0];
  _RAND_213 = {1{`RANDOM}};
  io_out_0_r_42_im = _RAND_213[16:0];
  _RAND_214 = {1{`RANDOM}};
  io_out_0_r_43_re = _RAND_214[16:0];
  _RAND_215 = {1{`RANDOM}};
  io_out_0_r_43_im = _RAND_215[16:0];
  _RAND_216 = {1{`RANDOM}};
  io_out_0_r_44_re = _RAND_216[16:0];
  _RAND_217 = {1{`RANDOM}};
  io_out_0_r_44_im = _RAND_217[16:0];
  _RAND_218 = {1{`RANDOM}};
  io_out_0_r_45_re = _RAND_218[16:0];
  _RAND_219 = {1{`RANDOM}};
  io_out_0_r_45_im = _RAND_219[16:0];
  _RAND_220 = {1{`RANDOM}};
  io_out_0_r_46_re = _RAND_220[16:0];
  _RAND_221 = {1{`RANDOM}};
  io_out_0_r_46_im = _RAND_221[16:0];
  _RAND_222 = {1{`RANDOM}};
  io_out_0_r_47_re = _RAND_222[16:0];
  _RAND_223 = {1{`RANDOM}};
  io_out_0_r_47_im = _RAND_223[16:0];
  _RAND_224 = {1{`RANDOM}};
  io_out_0_r_48_re = _RAND_224[16:0];
  _RAND_225 = {1{`RANDOM}};
  io_out_0_r_48_im = _RAND_225[16:0];
  _RAND_226 = {1{`RANDOM}};
  io_out_0_r_49_re = _RAND_226[16:0];
  _RAND_227 = {1{`RANDOM}};
  io_out_0_r_49_im = _RAND_227[16:0];
  _RAND_228 = {1{`RANDOM}};
  io_out_0_r_50_re = _RAND_228[16:0];
  _RAND_229 = {1{`RANDOM}};
  io_out_0_r_50_im = _RAND_229[16:0];
  _RAND_230 = {1{`RANDOM}};
  io_out_0_r_51_re = _RAND_230[16:0];
  _RAND_231 = {1{`RANDOM}};
  io_out_0_r_51_im = _RAND_231[16:0];
  _RAND_232 = {1{`RANDOM}};
  io_out_0_r_52_re = _RAND_232[16:0];
  _RAND_233 = {1{`RANDOM}};
  io_out_0_r_52_im = _RAND_233[16:0];
  _RAND_234 = {1{`RANDOM}};
  io_out_0_r_53_re = _RAND_234[16:0];
  _RAND_235 = {1{`RANDOM}};
  io_out_0_r_53_im = _RAND_235[16:0];
  _RAND_236 = {1{`RANDOM}};
  io_out_0_r_54_re = _RAND_236[16:0];
  _RAND_237 = {1{`RANDOM}};
  io_out_0_r_54_im = _RAND_237[16:0];
  _RAND_238 = {1{`RANDOM}};
  io_out_0_r_55_re = _RAND_238[16:0];
  _RAND_239 = {1{`RANDOM}};
  io_out_0_r_55_im = _RAND_239[16:0];
  _RAND_240 = {1{`RANDOM}};
  io_out_0_r_56_re = _RAND_240[16:0];
  _RAND_241 = {1{`RANDOM}};
  io_out_0_r_56_im = _RAND_241[16:0];
  _RAND_242 = {1{`RANDOM}};
  io_out_0_r_57_re = _RAND_242[16:0];
  _RAND_243 = {1{`RANDOM}};
  io_out_0_r_57_im = _RAND_243[16:0];
  _RAND_244 = {1{`RANDOM}};
  io_out_0_r_58_re = _RAND_244[16:0];
  _RAND_245 = {1{`RANDOM}};
  io_out_0_r_58_im = _RAND_245[16:0];
  _RAND_246 = {1{`RANDOM}};
  io_out_0_r_59_re = _RAND_246[16:0];
  _RAND_247 = {1{`RANDOM}};
  io_out_0_r_59_im = _RAND_247[16:0];
  _RAND_248 = {1{`RANDOM}};
  io_out_0_r_60_re = _RAND_248[16:0];
  _RAND_249 = {1{`RANDOM}};
  io_out_0_r_60_im = _RAND_249[16:0];
  _RAND_250 = {1{`RANDOM}};
  io_out_0_r_61_re = _RAND_250[16:0];
  _RAND_251 = {1{`RANDOM}};
  io_out_0_r_61_im = _RAND_251[16:0];
  _RAND_252 = {1{`RANDOM}};
  io_out_0_r_62_re = _RAND_252[16:0];
  _RAND_253 = {1{`RANDOM}};
  io_out_0_r_62_im = _RAND_253[16:0];
  _RAND_254 = {1{`RANDOM}};
  io_out_0_r_63_re = _RAND_254[16:0];
  _RAND_255 = {1{`RANDOM}};
  io_out_0_r_63_im = _RAND_255[16:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module Switch_1(
  input         clock,
  input  [16:0] io_in_0_re,
  input  [16:0] io_in_0_im,
  input  [16:0] io_in_1_re,
  input  [16:0] io_in_1_im,
  output [16:0] io_out_0_re,
  output [16:0] io_out_0_im,
  output [16:0] io_out_1_re,
  output [16:0] io_out_1_im,
  input         io_sel
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_9;
  reg [31:0] _RAND_10;
  reg [31:0] _RAND_11;
  reg [31:0] _RAND_12;
  reg [31:0] _RAND_13;
  reg [31:0] _RAND_14;
  reg [31:0] _RAND_15;
  reg [31:0] _RAND_16;
  reg [31:0] _RAND_17;
  reg [31:0] _RAND_18;
  reg [31:0] _RAND_19;
  reg [31:0] _RAND_20;
  reg [31:0] _RAND_21;
  reg [31:0] _RAND_22;
  reg [31:0] _RAND_23;
  reg [31:0] _RAND_24;
  reg [31:0] _RAND_25;
  reg [31:0] _RAND_26;
  reg [31:0] _RAND_27;
  reg [31:0] _RAND_28;
  reg [31:0] _RAND_29;
  reg [31:0] _RAND_30;
  reg [31:0] _RAND_31;
  reg [31:0] _RAND_32;
  reg [31:0] _RAND_33;
  reg [31:0] _RAND_34;
  reg [31:0] _RAND_35;
  reg [31:0] _RAND_36;
  reg [31:0] _RAND_37;
  reg [31:0] _RAND_38;
  reg [31:0] _RAND_39;
  reg [31:0] _RAND_40;
  reg [31:0] _RAND_41;
  reg [31:0] _RAND_42;
  reg [31:0] _RAND_43;
  reg [31:0] _RAND_44;
  reg [31:0] _RAND_45;
  reg [31:0] _RAND_46;
  reg [31:0] _RAND_47;
  reg [31:0] _RAND_48;
  reg [31:0] _RAND_49;
  reg [31:0] _RAND_50;
  reg [31:0] _RAND_51;
  reg [31:0] _RAND_52;
  reg [31:0] _RAND_53;
  reg [31:0] _RAND_54;
  reg [31:0] _RAND_55;
  reg [31:0] _RAND_56;
  reg [31:0] _RAND_57;
  reg [31:0] _RAND_58;
  reg [31:0] _RAND_59;
  reg [31:0] _RAND_60;
  reg [31:0] _RAND_61;
  reg [31:0] _RAND_62;
  reg [31:0] _RAND_63;
  reg [31:0] _RAND_64;
  reg [31:0] _RAND_65;
  reg [31:0] _RAND_66;
  reg [31:0] _RAND_67;
  reg [31:0] _RAND_68;
  reg [31:0] _RAND_69;
  reg [31:0] _RAND_70;
  reg [31:0] _RAND_71;
  reg [31:0] _RAND_72;
  reg [31:0] _RAND_73;
  reg [31:0] _RAND_74;
  reg [31:0] _RAND_75;
  reg [31:0] _RAND_76;
  reg [31:0] _RAND_77;
  reg [31:0] _RAND_78;
  reg [31:0] _RAND_79;
  reg [31:0] _RAND_80;
  reg [31:0] _RAND_81;
  reg [31:0] _RAND_82;
  reg [31:0] _RAND_83;
  reg [31:0] _RAND_84;
  reg [31:0] _RAND_85;
  reg [31:0] _RAND_86;
  reg [31:0] _RAND_87;
  reg [31:0] _RAND_88;
  reg [31:0] _RAND_89;
  reg [31:0] _RAND_90;
  reg [31:0] _RAND_91;
  reg [31:0] _RAND_92;
  reg [31:0] _RAND_93;
  reg [31:0] _RAND_94;
  reg [31:0] _RAND_95;
  reg [31:0] _RAND_96;
  reg [31:0] _RAND_97;
  reg [31:0] _RAND_98;
  reg [31:0] _RAND_99;
  reg [31:0] _RAND_100;
  reg [31:0] _RAND_101;
  reg [31:0] _RAND_102;
  reg [31:0] _RAND_103;
  reg [31:0] _RAND_104;
  reg [31:0] _RAND_105;
  reg [31:0] _RAND_106;
  reg [31:0] _RAND_107;
  reg [31:0] _RAND_108;
  reg [31:0] _RAND_109;
  reg [31:0] _RAND_110;
  reg [31:0] _RAND_111;
  reg [31:0] _RAND_112;
  reg [31:0] _RAND_113;
  reg [31:0] _RAND_114;
  reg [31:0] _RAND_115;
  reg [31:0] _RAND_116;
  reg [31:0] _RAND_117;
  reg [31:0] _RAND_118;
  reg [31:0] _RAND_119;
  reg [31:0] _RAND_120;
  reg [31:0] _RAND_121;
  reg [31:0] _RAND_122;
  reg [31:0] _RAND_123;
  reg [31:0] _RAND_124;
  reg [31:0] _RAND_125;
  reg [31:0] _RAND_126;
  reg [31:0] _RAND_127;
`endif // RANDOMIZE_REG_INIT
  reg [16:0] swdata_1_r_re; // @[Reg.scala 19:16]
  reg [16:0] swdata_1_r_im; // @[Reg.scala 19:16]
  reg [16:0] swdata_1_r_1_re; // @[Reg.scala 19:16]
  reg [16:0] swdata_1_r_1_im; // @[Reg.scala 19:16]
  reg [16:0] swdata_1_r_2_re; // @[Reg.scala 19:16]
  reg [16:0] swdata_1_r_2_im; // @[Reg.scala 19:16]
  reg [16:0] swdata_1_r_3_re; // @[Reg.scala 19:16]
  reg [16:0] swdata_1_r_3_im; // @[Reg.scala 19:16]
  reg [16:0] swdata_1_r_4_re; // @[Reg.scala 19:16]
  reg [16:0] swdata_1_r_4_im; // @[Reg.scala 19:16]
  reg [16:0] swdata_1_r_5_re; // @[Reg.scala 19:16]
  reg [16:0] swdata_1_r_5_im; // @[Reg.scala 19:16]
  reg [16:0] swdata_1_r_6_re; // @[Reg.scala 19:16]
  reg [16:0] swdata_1_r_6_im; // @[Reg.scala 19:16]
  reg [16:0] swdata_1_r_7_re; // @[Reg.scala 19:16]
  reg [16:0] swdata_1_r_7_im; // @[Reg.scala 19:16]
  reg [16:0] swdata_1_r_8_re; // @[Reg.scala 19:16]
  reg [16:0] swdata_1_r_8_im; // @[Reg.scala 19:16]
  reg [16:0] swdata_1_r_9_re; // @[Reg.scala 19:16]
  reg [16:0] swdata_1_r_9_im; // @[Reg.scala 19:16]
  reg [16:0] swdata_1_r_10_re; // @[Reg.scala 19:16]
  reg [16:0] swdata_1_r_10_im; // @[Reg.scala 19:16]
  reg [16:0] swdata_1_r_11_re; // @[Reg.scala 19:16]
  reg [16:0] swdata_1_r_11_im; // @[Reg.scala 19:16]
  reg [16:0] swdata_1_r_12_re; // @[Reg.scala 19:16]
  reg [16:0] swdata_1_r_12_im; // @[Reg.scala 19:16]
  reg [16:0] swdata_1_r_13_re; // @[Reg.scala 19:16]
  reg [16:0] swdata_1_r_13_im; // @[Reg.scala 19:16]
  reg [16:0] swdata_1_r_14_re; // @[Reg.scala 19:16]
  reg [16:0] swdata_1_r_14_im; // @[Reg.scala 19:16]
  reg [16:0] swdata_1_r_15_re; // @[Reg.scala 19:16]
  reg [16:0] swdata_1_r_15_im; // @[Reg.scala 19:16]
  reg [16:0] swdata_1_r_16_re; // @[Reg.scala 19:16]
  reg [16:0] swdata_1_r_16_im; // @[Reg.scala 19:16]
  reg [16:0] swdata_1_r_17_re; // @[Reg.scala 19:16]
  reg [16:0] swdata_1_r_17_im; // @[Reg.scala 19:16]
  reg [16:0] swdata_1_r_18_re; // @[Reg.scala 19:16]
  reg [16:0] swdata_1_r_18_im; // @[Reg.scala 19:16]
  reg [16:0] swdata_1_r_19_re; // @[Reg.scala 19:16]
  reg [16:0] swdata_1_r_19_im; // @[Reg.scala 19:16]
  reg [16:0] swdata_1_r_20_re; // @[Reg.scala 19:16]
  reg [16:0] swdata_1_r_20_im; // @[Reg.scala 19:16]
  reg [16:0] swdata_1_r_21_re; // @[Reg.scala 19:16]
  reg [16:0] swdata_1_r_21_im; // @[Reg.scala 19:16]
  reg [16:0] swdata_1_r_22_re; // @[Reg.scala 19:16]
  reg [16:0] swdata_1_r_22_im; // @[Reg.scala 19:16]
  reg [16:0] swdata_1_r_23_re; // @[Reg.scala 19:16]
  reg [16:0] swdata_1_r_23_im; // @[Reg.scala 19:16]
  reg [16:0] swdata_1_r_24_re; // @[Reg.scala 19:16]
  reg [16:0] swdata_1_r_24_im; // @[Reg.scala 19:16]
  reg [16:0] swdata_1_r_25_re; // @[Reg.scala 19:16]
  reg [16:0] swdata_1_r_25_im; // @[Reg.scala 19:16]
  reg [16:0] swdata_1_r_26_re; // @[Reg.scala 19:16]
  reg [16:0] swdata_1_r_26_im; // @[Reg.scala 19:16]
  reg [16:0] swdata_1_r_27_re; // @[Reg.scala 19:16]
  reg [16:0] swdata_1_r_27_im; // @[Reg.scala 19:16]
  reg [16:0] swdata_1_r_28_re; // @[Reg.scala 19:16]
  reg [16:0] swdata_1_r_28_im; // @[Reg.scala 19:16]
  reg [16:0] swdata_1_r_29_re; // @[Reg.scala 19:16]
  reg [16:0] swdata_1_r_29_im; // @[Reg.scala 19:16]
  reg [16:0] swdata_1_r_30_re; // @[Reg.scala 19:16]
  reg [16:0] swdata_1_r_30_im; // @[Reg.scala 19:16]
  reg [16:0] swdata_1_r_31_re; // @[Reg.scala 19:16]
  reg [16:0] swdata_1_r_31_im; // @[Reg.scala 19:16]
  reg [16:0] io_out_0_r_re; // @[Reg.scala 19:16]
  reg [16:0] io_out_0_r_im; // @[Reg.scala 19:16]
  reg [16:0] io_out_0_r_1_re; // @[Reg.scala 19:16]
  reg [16:0] io_out_0_r_1_im; // @[Reg.scala 19:16]
  reg [16:0] io_out_0_r_2_re; // @[Reg.scala 19:16]
  reg [16:0] io_out_0_r_2_im; // @[Reg.scala 19:16]
  reg [16:0] io_out_0_r_3_re; // @[Reg.scala 19:16]
  reg [16:0] io_out_0_r_3_im; // @[Reg.scala 19:16]
  reg [16:0] io_out_0_r_4_re; // @[Reg.scala 19:16]
  reg [16:0] io_out_0_r_4_im; // @[Reg.scala 19:16]
  reg [16:0] io_out_0_r_5_re; // @[Reg.scala 19:16]
  reg [16:0] io_out_0_r_5_im; // @[Reg.scala 19:16]
  reg [16:0] io_out_0_r_6_re; // @[Reg.scala 19:16]
  reg [16:0] io_out_0_r_6_im; // @[Reg.scala 19:16]
  reg [16:0] io_out_0_r_7_re; // @[Reg.scala 19:16]
  reg [16:0] io_out_0_r_7_im; // @[Reg.scala 19:16]
  reg [16:0] io_out_0_r_8_re; // @[Reg.scala 19:16]
  reg [16:0] io_out_0_r_8_im; // @[Reg.scala 19:16]
  reg [16:0] io_out_0_r_9_re; // @[Reg.scala 19:16]
  reg [16:0] io_out_0_r_9_im; // @[Reg.scala 19:16]
  reg [16:0] io_out_0_r_10_re; // @[Reg.scala 19:16]
  reg [16:0] io_out_0_r_10_im; // @[Reg.scala 19:16]
  reg [16:0] io_out_0_r_11_re; // @[Reg.scala 19:16]
  reg [16:0] io_out_0_r_11_im; // @[Reg.scala 19:16]
  reg [16:0] io_out_0_r_12_re; // @[Reg.scala 19:16]
  reg [16:0] io_out_0_r_12_im; // @[Reg.scala 19:16]
  reg [16:0] io_out_0_r_13_re; // @[Reg.scala 19:16]
  reg [16:0] io_out_0_r_13_im; // @[Reg.scala 19:16]
  reg [16:0] io_out_0_r_14_re; // @[Reg.scala 19:16]
  reg [16:0] io_out_0_r_14_im; // @[Reg.scala 19:16]
  reg [16:0] io_out_0_r_15_re; // @[Reg.scala 19:16]
  reg [16:0] io_out_0_r_15_im; // @[Reg.scala 19:16]
  reg [16:0] io_out_0_r_16_re; // @[Reg.scala 19:16]
  reg [16:0] io_out_0_r_16_im; // @[Reg.scala 19:16]
  reg [16:0] io_out_0_r_17_re; // @[Reg.scala 19:16]
  reg [16:0] io_out_0_r_17_im; // @[Reg.scala 19:16]
  reg [16:0] io_out_0_r_18_re; // @[Reg.scala 19:16]
  reg [16:0] io_out_0_r_18_im; // @[Reg.scala 19:16]
  reg [16:0] io_out_0_r_19_re; // @[Reg.scala 19:16]
  reg [16:0] io_out_0_r_19_im; // @[Reg.scala 19:16]
  reg [16:0] io_out_0_r_20_re; // @[Reg.scala 19:16]
  reg [16:0] io_out_0_r_20_im; // @[Reg.scala 19:16]
  reg [16:0] io_out_0_r_21_re; // @[Reg.scala 19:16]
  reg [16:0] io_out_0_r_21_im; // @[Reg.scala 19:16]
  reg [16:0] io_out_0_r_22_re; // @[Reg.scala 19:16]
  reg [16:0] io_out_0_r_22_im; // @[Reg.scala 19:16]
  reg [16:0] io_out_0_r_23_re; // @[Reg.scala 19:16]
  reg [16:0] io_out_0_r_23_im; // @[Reg.scala 19:16]
  reg [16:0] io_out_0_r_24_re; // @[Reg.scala 19:16]
  reg [16:0] io_out_0_r_24_im; // @[Reg.scala 19:16]
  reg [16:0] io_out_0_r_25_re; // @[Reg.scala 19:16]
  reg [16:0] io_out_0_r_25_im; // @[Reg.scala 19:16]
  reg [16:0] io_out_0_r_26_re; // @[Reg.scala 19:16]
  reg [16:0] io_out_0_r_26_im; // @[Reg.scala 19:16]
  reg [16:0] io_out_0_r_27_re; // @[Reg.scala 19:16]
  reg [16:0] io_out_0_r_27_im; // @[Reg.scala 19:16]
  reg [16:0] io_out_0_r_28_re; // @[Reg.scala 19:16]
  reg [16:0] io_out_0_r_28_im; // @[Reg.scala 19:16]
  reg [16:0] io_out_0_r_29_re; // @[Reg.scala 19:16]
  reg [16:0] io_out_0_r_29_im; // @[Reg.scala 19:16]
  reg [16:0] io_out_0_r_30_re; // @[Reg.scala 19:16]
  reg [16:0] io_out_0_r_30_im; // @[Reg.scala 19:16]
  reg [16:0] io_out_0_r_31_re; // @[Reg.scala 19:16]
  reg [16:0] io_out_0_r_31_im; // @[Reg.scala 19:16]
  assign io_out_0_re = io_out_0_r_31_re; // @[Modules.scala 306:38]
  assign io_out_0_im = io_out_0_r_31_im; // @[Modules.scala 306:38]
  assign io_out_1_re = io_sel ? io_in_0_re : swdata_1_r_31_re; // @[Modules.scala 306:{38,38}]
  assign io_out_1_im = io_sel ? io_in_0_im : swdata_1_r_31_im; // @[Modules.scala 306:{38,38}]
  always @(posedge clock) begin
    swdata_1_r_re <= io_in_1_re; // @[Reg.scala 19:16 20:{18,22}]
    swdata_1_r_im <= io_in_1_im; // @[Reg.scala 19:16 20:{18,22}]
    swdata_1_r_1_re <= swdata_1_r_re; // @[Reg.scala 19:16 20:{18,22}]
    swdata_1_r_1_im <= swdata_1_r_im; // @[Reg.scala 19:16 20:{18,22}]
    swdata_1_r_2_re <= swdata_1_r_1_re; // @[Reg.scala 19:16 20:{18,22}]
    swdata_1_r_2_im <= swdata_1_r_1_im; // @[Reg.scala 19:16 20:{18,22}]
    swdata_1_r_3_re <= swdata_1_r_2_re; // @[Reg.scala 19:16 20:{18,22}]
    swdata_1_r_3_im <= swdata_1_r_2_im; // @[Reg.scala 19:16 20:{18,22}]
    swdata_1_r_4_re <= swdata_1_r_3_re; // @[Reg.scala 19:16 20:{18,22}]
    swdata_1_r_4_im <= swdata_1_r_3_im; // @[Reg.scala 19:16 20:{18,22}]
    swdata_1_r_5_re <= swdata_1_r_4_re; // @[Reg.scala 19:16 20:{18,22}]
    swdata_1_r_5_im <= swdata_1_r_4_im; // @[Reg.scala 19:16 20:{18,22}]
    swdata_1_r_6_re <= swdata_1_r_5_re; // @[Reg.scala 19:16 20:{18,22}]
    swdata_1_r_6_im <= swdata_1_r_5_im; // @[Reg.scala 19:16 20:{18,22}]
    swdata_1_r_7_re <= swdata_1_r_6_re; // @[Reg.scala 19:16 20:{18,22}]
    swdata_1_r_7_im <= swdata_1_r_6_im; // @[Reg.scala 19:16 20:{18,22}]
    swdata_1_r_8_re <= swdata_1_r_7_re; // @[Reg.scala 19:16 20:{18,22}]
    swdata_1_r_8_im <= swdata_1_r_7_im; // @[Reg.scala 19:16 20:{18,22}]
    swdata_1_r_9_re <= swdata_1_r_8_re; // @[Reg.scala 19:16 20:{18,22}]
    swdata_1_r_9_im <= swdata_1_r_8_im; // @[Reg.scala 19:16 20:{18,22}]
    swdata_1_r_10_re <= swdata_1_r_9_re; // @[Reg.scala 19:16 20:{18,22}]
    swdata_1_r_10_im <= swdata_1_r_9_im; // @[Reg.scala 19:16 20:{18,22}]
    swdata_1_r_11_re <= swdata_1_r_10_re; // @[Reg.scala 19:16 20:{18,22}]
    swdata_1_r_11_im <= swdata_1_r_10_im; // @[Reg.scala 19:16 20:{18,22}]
    swdata_1_r_12_re <= swdata_1_r_11_re; // @[Reg.scala 19:16 20:{18,22}]
    swdata_1_r_12_im <= swdata_1_r_11_im; // @[Reg.scala 19:16 20:{18,22}]
    swdata_1_r_13_re <= swdata_1_r_12_re; // @[Reg.scala 19:16 20:{18,22}]
    swdata_1_r_13_im <= swdata_1_r_12_im; // @[Reg.scala 19:16 20:{18,22}]
    swdata_1_r_14_re <= swdata_1_r_13_re; // @[Reg.scala 19:16 20:{18,22}]
    swdata_1_r_14_im <= swdata_1_r_13_im; // @[Reg.scala 19:16 20:{18,22}]
    swdata_1_r_15_re <= swdata_1_r_14_re; // @[Reg.scala 19:16 20:{18,22}]
    swdata_1_r_15_im <= swdata_1_r_14_im; // @[Reg.scala 19:16 20:{18,22}]
    swdata_1_r_16_re <= swdata_1_r_15_re; // @[Reg.scala 19:16 20:{18,22}]
    swdata_1_r_16_im <= swdata_1_r_15_im; // @[Reg.scala 19:16 20:{18,22}]
    swdata_1_r_17_re <= swdata_1_r_16_re; // @[Reg.scala 19:16 20:{18,22}]
    swdata_1_r_17_im <= swdata_1_r_16_im; // @[Reg.scala 19:16 20:{18,22}]
    swdata_1_r_18_re <= swdata_1_r_17_re; // @[Reg.scala 19:16 20:{18,22}]
    swdata_1_r_18_im <= swdata_1_r_17_im; // @[Reg.scala 19:16 20:{18,22}]
    swdata_1_r_19_re <= swdata_1_r_18_re; // @[Reg.scala 19:16 20:{18,22}]
    swdata_1_r_19_im <= swdata_1_r_18_im; // @[Reg.scala 19:16 20:{18,22}]
    swdata_1_r_20_re <= swdata_1_r_19_re; // @[Reg.scala 19:16 20:{18,22}]
    swdata_1_r_20_im <= swdata_1_r_19_im; // @[Reg.scala 19:16 20:{18,22}]
    swdata_1_r_21_re <= swdata_1_r_20_re; // @[Reg.scala 19:16 20:{18,22}]
    swdata_1_r_21_im <= swdata_1_r_20_im; // @[Reg.scala 19:16 20:{18,22}]
    swdata_1_r_22_re <= swdata_1_r_21_re; // @[Reg.scala 19:16 20:{18,22}]
    swdata_1_r_22_im <= swdata_1_r_21_im; // @[Reg.scala 19:16 20:{18,22}]
    swdata_1_r_23_re <= swdata_1_r_22_re; // @[Reg.scala 19:16 20:{18,22}]
    swdata_1_r_23_im <= swdata_1_r_22_im; // @[Reg.scala 19:16 20:{18,22}]
    swdata_1_r_24_re <= swdata_1_r_23_re; // @[Reg.scala 19:16 20:{18,22}]
    swdata_1_r_24_im <= swdata_1_r_23_im; // @[Reg.scala 19:16 20:{18,22}]
    swdata_1_r_25_re <= swdata_1_r_24_re; // @[Reg.scala 19:16 20:{18,22}]
    swdata_1_r_25_im <= swdata_1_r_24_im; // @[Reg.scala 19:16 20:{18,22}]
    swdata_1_r_26_re <= swdata_1_r_25_re; // @[Reg.scala 19:16 20:{18,22}]
    swdata_1_r_26_im <= swdata_1_r_25_im; // @[Reg.scala 19:16 20:{18,22}]
    swdata_1_r_27_re <= swdata_1_r_26_re; // @[Reg.scala 19:16 20:{18,22}]
    swdata_1_r_27_im <= swdata_1_r_26_im; // @[Reg.scala 19:16 20:{18,22}]
    swdata_1_r_28_re <= swdata_1_r_27_re; // @[Reg.scala 19:16 20:{18,22}]
    swdata_1_r_28_im <= swdata_1_r_27_im; // @[Reg.scala 19:16 20:{18,22}]
    swdata_1_r_29_re <= swdata_1_r_28_re; // @[Reg.scala 19:16 20:{18,22}]
    swdata_1_r_29_im <= swdata_1_r_28_im; // @[Reg.scala 19:16 20:{18,22}]
    swdata_1_r_30_re <= swdata_1_r_29_re; // @[Reg.scala 19:16 20:{18,22}]
    swdata_1_r_30_im <= swdata_1_r_29_im; // @[Reg.scala 19:16 20:{18,22}]
    swdata_1_r_31_re <= swdata_1_r_30_re; // @[Reg.scala 19:16 20:{18,22}]
    swdata_1_r_31_im <= swdata_1_r_30_im; // @[Reg.scala 19:16 20:{18,22}]
    if (io_sel) begin // @[Reg.scala 20:22]
      io_out_0_r_re <= swdata_1_r_31_re; // @[Reg.scala 20:22]
    end else begin
      io_out_0_r_re <= io_in_0_re;
    end
    if (io_sel) begin // @[Reg.scala 20:22]
      io_out_0_r_im <= swdata_1_r_31_im; // @[Reg.scala 20:22]
    end else begin
      io_out_0_r_im <= io_in_0_im;
    end
    io_out_0_r_1_re <= io_out_0_r_re; // @[Reg.scala 19:16 20:{18,22}]
    io_out_0_r_1_im <= io_out_0_r_im; // @[Reg.scala 19:16 20:{18,22}]
    io_out_0_r_2_re <= io_out_0_r_1_re; // @[Reg.scala 19:16 20:{18,22}]
    io_out_0_r_2_im <= io_out_0_r_1_im; // @[Reg.scala 19:16 20:{18,22}]
    io_out_0_r_3_re <= io_out_0_r_2_re; // @[Reg.scala 19:16 20:{18,22}]
    io_out_0_r_3_im <= io_out_0_r_2_im; // @[Reg.scala 19:16 20:{18,22}]
    io_out_0_r_4_re <= io_out_0_r_3_re; // @[Reg.scala 19:16 20:{18,22}]
    io_out_0_r_4_im <= io_out_0_r_3_im; // @[Reg.scala 19:16 20:{18,22}]
    io_out_0_r_5_re <= io_out_0_r_4_re; // @[Reg.scala 19:16 20:{18,22}]
    io_out_0_r_5_im <= io_out_0_r_4_im; // @[Reg.scala 19:16 20:{18,22}]
    io_out_0_r_6_re <= io_out_0_r_5_re; // @[Reg.scala 19:16 20:{18,22}]
    io_out_0_r_6_im <= io_out_0_r_5_im; // @[Reg.scala 19:16 20:{18,22}]
    io_out_0_r_7_re <= io_out_0_r_6_re; // @[Reg.scala 19:16 20:{18,22}]
    io_out_0_r_7_im <= io_out_0_r_6_im; // @[Reg.scala 19:16 20:{18,22}]
    io_out_0_r_8_re <= io_out_0_r_7_re; // @[Reg.scala 19:16 20:{18,22}]
    io_out_0_r_8_im <= io_out_0_r_7_im; // @[Reg.scala 19:16 20:{18,22}]
    io_out_0_r_9_re <= io_out_0_r_8_re; // @[Reg.scala 19:16 20:{18,22}]
    io_out_0_r_9_im <= io_out_0_r_8_im; // @[Reg.scala 19:16 20:{18,22}]
    io_out_0_r_10_re <= io_out_0_r_9_re; // @[Reg.scala 19:16 20:{18,22}]
    io_out_0_r_10_im <= io_out_0_r_9_im; // @[Reg.scala 19:16 20:{18,22}]
    io_out_0_r_11_re <= io_out_0_r_10_re; // @[Reg.scala 19:16 20:{18,22}]
    io_out_0_r_11_im <= io_out_0_r_10_im; // @[Reg.scala 19:16 20:{18,22}]
    io_out_0_r_12_re <= io_out_0_r_11_re; // @[Reg.scala 19:16 20:{18,22}]
    io_out_0_r_12_im <= io_out_0_r_11_im; // @[Reg.scala 19:16 20:{18,22}]
    io_out_0_r_13_re <= io_out_0_r_12_re; // @[Reg.scala 19:16 20:{18,22}]
    io_out_0_r_13_im <= io_out_0_r_12_im; // @[Reg.scala 19:16 20:{18,22}]
    io_out_0_r_14_re <= io_out_0_r_13_re; // @[Reg.scala 19:16 20:{18,22}]
    io_out_0_r_14_im <= io_out_0_r_13_im; // @[Reg.scala 19:16 20:{18,22}]
    io_out_0_r_15_re <= io_out_0_r_14_re; // @[Reg.scala 19:16 20:{18,22}]
    io_out_0_r_15_im <= io_out_0_r_14_im; // @[Reg.scala 19:16 20:{18,22}]
    io_out_0_r_16_re <= io_out_0_r_15_re; // @[Reg.scala 19:16 20:{18,22}]
    io_out_0_r_16_im <= io_out_0_r_15_im; // @[Reg.scala 19:16 20:{18,22}]
    io_out_0_r_17_re <= io_out_0_r_16_re; // @[Reg.scala 19:16 20:{18,22}]
    io_out_0_r_17_im <= io_out_0_r_16_im; // @[Reg.scala 19:16 20:{18,22}]
    io_out_0_r_18_re <= io_out_0_r_17_re; // @[Reg.scala 19:16 20:{18,22}]
    io_out_0_r_18_im <= io_out_0_r_17_im; // @[Reg.scala 19:16 20:{18,22}]
    io_out_0_r_19_re <= io_out_0_r_18_re; // @[Reg.scala 19:16 20:{18,22}]
    io_out_0_r_19_im <= io_out_0_r_18_im; // @[Reg.scala 19:16 20:{18,22}]
    io_out_0_r_20_re <= io_out_0_r_19_re; // @[Reg.scala 19:16 20:{18,22}]
    io_out_0_r_20_im <= io_out_0_r_19_im; // @[Reg.scala 19:16 20:{18,22}]
    io_out_0_r_21_re <= io_out_0_r_20_re; // @[Reg.scala 19:16 20:{18,22}]
    io_out_0_r_21_im <= io_out_0_r_20_im; // @[Reg.scala 19:16 20:{18,22}]
    io_out_0_r_22_re <= io_out_0_r_21_re; // @[Reg.scala 19:16 20:{18,22}]
    io_out_0_r_22_im <= io_out_0_r_21_im; // @[Reg.scala 19:16 20:{18,22}]
    io_out_0_r_23_re <= io_out_0_r_22_re; // @[Reg.scala 19:16 20:{18,22}]
    io_out_0_r_23_im <= io_out_0_r_22_im; // @[Reg.scala 19:16 20:{18,22}]
    io_out_0_r_24_re <= io_out_0_r_23_re; // @[Reg.scala 19:16 20:{18,22}]
    io_out_0_r_24_im <= io_out_0_r_23_im; // @[Reg.scala 19:16 20:{18,22}]
    io_out_0_r_25_re <= io_out_0_r_24_re; // @[Reg.scala 19:16 20:{18,22}]
    io_out_0_r_25_im <= io_out_0_r_24_im; // @[Reg.scala 19:16 20:{18,22}]
    io_out_0_r_26_re <= io_out_0_r_25_re; // @[Reg.scala 19:16 20:{18,22}]
    io_out_0_r_26_im <= io_out_0_r_25_im; // @[Reg.scala 19:16 20:{18,22}]
    io_out_0_r_27_re <= io_out_0_r_26_re; // @[Reg.scala 19:16 20:{18,22}]
    io_out_0_r_27_im <= io_out_0_r_26_im; // @[Reg.scala 19:16 20:{18,22}]
    io_out_0_r_28_re <= io_out_0_r_27_re; // @[Reg.scala 19:16 20:{18,22}]
    io_out_0_r_28_im <= io_out_0_r_27_im; // @[Reg.scala 19:16 20:{18,22}]
    io_out_0_r_29_re <= io_out_0_r_28_re; // @[Reg.scala 19:16 20:{18,22}]
    io_out_0_r_29_im <= io_out_0_r_28_im; // @[Reg.scala 19:16 20:{18,22}]
    io_out_0_r_30_re <= io_out_0_r_29_re; // @[Reg.scala 19:16 20:{18,22}]
    io_out_0_r_30_im <= io_out_0_r_29_im; // @[Reg.scala 19:16 20:{18,22}]
    io_out_0_r_31_re <= io_out_0_r_30_re; // @[Reg.scala 19:16 20:{18,22}]
    io_out_0_r_31_im <= io_out_0_r_30_im; // @[Reg.scala 19:16 20:{18,22}]
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  swdata_1_r_re = _RAND_0[16:0];
  _RAND_1 = {1{`RANDOM}};
  swdata_1_r_im = _RAND_1[16:0];
  _RAND_2 = {1{`RANDOM}};
  swdata_1_r_1_re = _RAND_2[16:0];
  _RAND_3 = {1{`RANDOM}};
  swdata_1_r_1_im = _RAND_3[16:0];
  _RAND_4 = {1{`RANDOM}};
  swdata_1_r_2_re = _RAND_4[16:0];
  _RAND_5 = {1{`RANDOM}};
  swdata_1_r_2_im = _RAND_5[16:0];
  _RAND_6 = {1{`RANDOM}};
  swdata_1_r_3_re = _RAND_6[16:0];
  _RAND_7 = {1{`RANDOM}};
  swdata_1_r_3_im = _RAND_7[16:0];
  _RAND_8 = {1{`RANDOM}};
  swdata_1_r_4_re = _RAND_8[16:0];
  _RAND_9 = {1{`RANDOM}};
  swdata_1_r_4_im = _RAND_9[16:0];
  _RAND_10 = {1{`RANDOM}};
  swdata_1_r_5_re = _RAND_10[16:0];
  _RAND_11 = {1{`RANDOM}};
  swdata_1_r_5_im = _RAND_11[16:0];
  _RAND_12 = {1{`RANDOM}};
  swdata_1_r_6_re = _RAND_12[16:0];
  _RAND_13 = {1{`RANDOM}};
  swdata_1_r_6_im = _RAND_13[16:0];
  _RAND_14 = {1{`RANDOM}};
  swdata_1_r_7_re = _RAND_14[16:0];
  _RAND_15 = {1{`RANDOM}};
  swdata_1_r_7_im = _RAND_15[16:0];
  _RAND_16 = {1{`RANDOM}};
  swdata_1_r_8_re = _RAND_16[16:0];
  _RAND_17 = {1{`RANDOM}};
  swdata_1_r_8_im = _RAND_17[16:0];
  _RAND_18 = {1{`RANDOM}};
  swdata_1_r_9_re = _RAND_18[16:0];
  _RAND_19 = {1{`RANDOM}};
  swdata_1_r_9_im = _RAND_19[16:0];
  _RAND_20 = {1{`RANDOM}};
  swdata_1_r_10_re = _RAND_20[16:0];
  _RAND_21 = {1{`RANDOM}};
  swdata_1_r_10_im = _RAND_21[16:0];
  _RAND_22 = {1{`RANDOM}};
  swdata_1_r_11_re = _RAND_22[16:0];
  _RAND_23 = {1{`RANDOM}};
  swdata_1_r_11_im = _RAND_23[16:0];
  _RAND_24 = {1{`RANDOM}};
  swdata_1_r_12_re = _RAND_24[16:0];
  _RAND_25 = {1{`RANDOM}};
  swdata_1_r_12_im = _RAND_25[16:0];
  _RAND_26 = {1{`RANDOM}};
  swdata_1_r_13_re = _RAND_26[16:0];
  _RAND_27 = {1{`RANDOM}};
  swdata_1_r_13_im = _RAND_27[16:0];
  _RAND_28 = {1{`RANDOM}};
  swdata_1_r_14_re = _RAND_28[16:0];
  _RAND_29 = {1{`RANDOM}};
  swdata_1_r_14_im = _RAND_29[16:0];
  _RAND_30 = {1{`RANDOM}};
  swdata_1_r_15_re = _RAND_30[16:0];
  _RAND_31 = {1{`RANDOM}};
  swdata_1_r_15_im = _RAND_31[16:0];
  _RAND_32 = {1{`RANDOM}};
  swdata_1_r_16_re = _RAND_32[16:0];
  _RAND_33 = {1{`RANDOM}};
  swdata_1_r_16_im = _RAND_33[16:0];
  _RAND_34 = {1{`RANDOM}};
  swdata_1_r_17_re = _RAND_34[16:0];
  _RAND_35 = {1{`RANDOM}};
  swdata_1_r_17_im = _RAND_35[16:0];
  _RAND_36 = {1{`RANDOM}};
  swdata_1_r_18_re = _RAND_36[16:0];
  _RAND_37 = {1{`RANDOM}};
  swdata_1_r_18_im = _RAND_37[16:0];
  _RAND_38 = {1{`RANDOM}};
  swdata_1_r_19_re = _RAND_38[16:0];
  _RAND_39 = {1{`RANDOM}};
  swdata_1_r_19_im = _RAND_39[16:0];
  _RAND_40 = {1{`RANDOM}};
  swdata_1_r_20_re = _RAND_40[16:0];
  _RAND_41 = {1{`RANDOM}};
  swdata_1_r_20_im = _RAND_41[16:0];
  _RAND_42 = {1{`RANDOM}};
  swdata_1_r_21_re = _RAND_42[16:0];
  _RAND_43 = {1{`RANDOM}};
  swdata_1_r_21_im = _RAND_43[16:0];
  _RAND_44 = {1{`RANDOM}};
  swdata_1_r_22_re = _RAND_44[16:0];
  _RAND_45 = {1{`RANDOM}};
  swdata_1_r_22_im = _RAND_45[16:0];
  _RAND_46 = {1{`RANDOM}};
  swdata_1_r_23_re = _RAND_46[16:0];
  _RAND_47 = {1{`RANDOM}};
  swdata_1_r_23_im = _RAND_47[16:0];
  _RAND_48 = {1{`RANDOM}};
  swdata_1_r_24_re = _RAND_48[16:0];
  _RAND_49 = {1{`RANDOM}};
  swdata_1_r_24_im = _RAND_49[16:0];
  _RAND_50 = {1{`RANDOM}};
  swdata_1_r_25_re = _RAND_50[16:0];
  _RAND_51 = {1{`RANDOM}};
  swdata_1_r_25_im = _RAND_51[16:0];
  _RAND_52 = {1{`RANDOM}};
  swdata_1_r_26_re = _RAND_52[16:0];
  _RAND_53 = {1{`RANDOM}};
  swdata_1_r_26_im = _RAND_53[16:0];
  _RAND_54 = {1{`RANDOM}};
  swdata_1_r_27_re = _RAND_54[16:0];
  _RAND_55 = {1{`RANDOM}};
  swdata_1_r_27_im = _RAND_55[16:0];
  _RAND_56 = {1{`RANDOM}};
  swdata_1_r_28_re = _RAND_56[16:0];
  _RAND_57 = {1{`RANDOM}};
  swdata_1_r_28_im = _RAND_57[16:0];
  _RAND_58 = {1{`RANDOM}};
  swdata_1_r_29_re = _RAND_58[16:0];
  _RAND_59 = {1{`RANDOM}};
  swdata_1_r_29_im = _RAND_59[16:0];
  _RAND_60 = {1{`RANDOM}};
  swdata_1_r_30_re = _RAND_60[16:0];
  _RAND_61 = {1{`RANDOM}};
  swdata_1_r_30_im = _RAND_61[16:0];
  _RAND_62 = {1{`RANDOM}};
  swdata_1_r_31_re = _RAND_62[16:0];
  _RAND_63 = {1{`RANDOM}};
  swdata_1_r_31_im = _RAND_63[16:0];
  _RAND_64 = {1{`RANDOM}};
  io_out_0_r_re = _RAND_64[16:0];
  _RAND_65 = {1{`RANDOM}};
  io_out_0_r_im = _RAND_65[16:0];
  _RAND_66 = {1{`RANDOM}};
  io_out_0_r_1_re = _RAND_66[16:0];
  _RAND_67 = {1{`RANDOM}};
  io_out_0_r_1_im = _RAND_67[16:0];
  _RAND_68 = {1{`RANDOM}};
  io_out_0_r_2_re = _RAND_68[16:0];
  _RAND_69 = {1{`RANDOM}};
  io_out_0_r_2_im = _RAND_69[16:0];
  _RAND_70 = {1{`RANDOM}};
  io_out_0_r_3_re = _RAND_70[16:0];
  _RAND_71 = {1{`RANDOM}};
  io_out_0_r_3_im = _RAND_71[16:0];
  _RAND_72 = {1{`RANDOM}};
  io_out_0_r_4_re = _RAND_72[16:0];
  _RAND_73 = {1{`RANDOM}};
  io_out_0_r_4_im = _RAND_73[16:0];
  _RAND_74 = {1{`RANDOM}};
  io_out_0_r_5_re = _RAND_74[16:0];
  _RAND_75 = {1{`RANDOM}};
  io_out_0_r_5_im = _RAND_75[16:0];
  _RAND_76 = {1{`RANDOM}};
  io_out_0_r_6_re = _RAND_76[16:0];
  _RAND_77 = {1{`RANDOM}};
  io_out_0_r_6_im = _RAND_77[16:0];
  _RAND_78 = {1{`RANDOM}};
  io_out_0_r_7_re = _RAND_78[16:0];
  _RAND_79 = {1{`RANDOM}};
  io_out_0_r_7_im = _RAND_79[16:0];
  _RAND_80 = {1{`RANDOM}};
  io_out_0_r_8_re = _RAND_80[16:0];
  _RAND_81 = {1{`RANDOM}};
  io_out_0_r_8_im = _RAND_81[16:0];
  _RAND_82 = {1{`RANDOM}};
  io_out_0_r_9_re = _RAND_82[16:0];
  _RAND_83 = {1{`RANDOM}};
  io_out_0_r_9_im = _RAND_83[16:0];
  _RAND_84 = {1{`RANDOM}};
  io_out_0_r_10_re = _RAND_84[16:0];
  _RAND_85 = {1{`RANDOM}};
  io_out_0_r_10_im = _RAND_85[16:0];
  _RAND_86 = {1{`RANDOM}};
  io_out_0_r_11_re = _RAND_86[16:0];
  _RAND_87 = {1{`RANDOM}};
  io_out_0_r_11_im = _RAND_87[16:0];
  _RAND_88 = {1{`RANDOM}};
  io_out_0_r_12_re = _RAND_88[16:0];
  _RAND_89 = {1{`RANDOM}};
  io_out_0_r_12_im = _RAND_89[16:0];
  _RAND_90 = {1{`RANDOM}};
  io_out_0_r_13_re = _RAND_90[16:0];
  _RAND_91 = {1{`RANDOM}};
  io_out_0_r_13_im = _RAND_91[16:0];
  _RAND_92 = {1{`RANDOM}};
  io_out_0_r_14_re = _RAND_92[16:0];
  _RAND_93 = {1{`RANDOM}};
  io_out_0_r_14_im = _RAND_93[16:0];
  _RAND_94 = {1{`RANDOM}};
  io_out_0_r_15_re = _RAND_94[16:0];
  _RAND_95 = {1{`RANDOM}};
  io_out_0_r_15_im = _RAND_95[16:0];
  _RAND_96 = {1{`RANDOM}};
  io_out_0_r_16_re = _RAND_96[16:0];
  _RAND_97 = {1{`RANDOM}};
  io_out_0_r_16_im = _RAND_97[16:0];
  _RAND_98 = {1{`RANDOM}};
  io_out_0_r_17_re = _RAND_98[16:0];
  _RAND_99 = {1{`RANDOM}};
  io_out_0_r_17_im = _RAND_99[16:0];
  _RAND_100 = {1{`RANDOM}};
  io_out_0_r_18_re = _RAND_100[16:0];
  _RAND_101 = {1{`RANDOM}};
  io_out_0_r_18_im = _RAND_101[16:0];
  _RAND_102 = {1{`RANDOM}};
  io_out_0_r_19_re = _RAND_102[16:0];
  _RAND_103 = {1{`RANDOM}};
  io_out_0_r_19_im = _RAND_103[16:0];
  _RAND_104 = {1{`RANDOM}};
  io_out_0_r_20_re = _RAND_104[16:0];
  _RAND_105 = {1{`RANDOM}};
  io_out_0_r_20_im = _RAND_105[16:0];
  _RAND_106 = {1{`RANDOM}};
  io_out_0_r_21_re = _RAND_106[16:0];
  _RAND_107 = {1{`RANDOM}};
  io_out_0_r_21_im = _RAND_107[16:0];
  _RAND_108 = {1{`RANDOM}};
  io_out_0_r_22_re = _RAND_108[16:0];
  _RAND_109 = {1{`RANDOM}};
  io_out_0_r_22_im = _RAND_109[16:0];
  _RAND_110 = {1{`RANDOM}};
  io_out_0_r_23_re = _RAND_110[16:0];
  _RAND_111 = {1{`RANDOM}};
  io_out_0_r_23_im = _RAND_111[16:0];
  _RAND_112 = {1{`RANDOM}};
  io_out_0_r_24_re = _RAND_112[16:0];
  _RAND_113 = {1{`RANDOM}};
  io_out_0_r_24_im = _RAND_113[16:0];
  _RAND_114 = {1{`RANDOM}};
  io_out_0_r_25_re = _RAND_114[16:0];
  _RAND_115 = {1{`RANDOM}};
  io_out_0_r_25_im = _RAND_115[16:0];
  _RAND_116 = {1{`RANDOM}};
  io_out_0_r_26_re = _RAND_116[16:0];
  _RAND_117 = {1{`RANDOM}};
  io_out_0_r_26_im = _RAND_117[16:0];
  _RAND_118 = {1{`RANDOM}};
  io_out_0_r_27_re = _RAND_118[16:0];
  _RAND_119 = {1{`RANDOM}};
  io_out_0_r_27_im = _RAND_119[16:0];
  _RAND_120 = {1{`RANDOM}};
  io_out_0_r_28_re = _RAND_120[16:0];
  _RAND_121 = {1{`RANDOM}};
  io_out_0_r_28_im = _RAND_121[16:0];
  _RAND_122 = {1{`RANDOM}};
  io_out_0_r_29_re = _RAND_122[16:0];
  _RAND_123 = {1{`RANDOM}};
  io_out_0_r_29_im = _RAND_123[16:0];
  _RAND_124 = {1{`RANDOM}};
  io_out_0_r_30_re = _RAND_124[16:0];
  _RAND_125 = {1{`RANDOM}};
  io_out_0_r_30_im = _RAND_125[16:0];
  _RAND_126 = {1{`RANDOM}};
  io_out_0_r_31_re = _RAND_126[16:0];
  _RAND_127 = {1{`RANDOM}};
  io_out_0_r_31_im = _RAND_127[16:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module Switch_2(
  input         clock,
  input  [16:0] io_in_0_re,
  input  [16:0] io_in_0_im,
  input  [16:0] io_in_1_re,
  input  [16:0] io_in_1_im,
  output [16:0] io_out_0_re,
  output [16:0] io_out_0_im,
  output [16:0] io_out_1_re,
  output [16:0] io_out_1_im,
  input         io_sel
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_9;
  reg [31:0] _RAND_10;
  reg [31:0] _RAND_11;
  reg [31:0] _RAND_12;
  reg [31:0] _RAND_13;
  reg [31:0] _RAND_14;
  reg [31:0] _RAND_15;
  reg [31:0] _RAND_16;
  reg [31:0] _RAND_17;
  reg [31:0] _RAND_18;
  reg [31:0] _RAND_19;
  reg [31:0] _RAND_20;
  reg [31:0] _RAND_21;
  reg [31:0] _RAND_22;
  reg [31:0] _RAND_23;
  reg [31:0] _RAND_24;
  reg [31:0] _RAND_25;
  reg [31:0] _RAND_26;
  reg [31:0] _RAND_27;
  reg [31:0] _RAND_28;
  reg [31:0] _RAND_29;
  reg [31:0] _RAND_30;
  reg [31:0] _RAND_31;
  reg [31:0] _RAND_32;
  reg [31:0] _RAND_33;
  reg [31:0] _RAND_34;
  reg [31:0] _RAND_35;
  reg [31:0] _RAND_36;
  reg [31:0] _RAND_37;
  reg [31:0] _RAND_38;
  reg [31:0] _RAND_39;
  reg [31:0] _RAND_40;
  reg [31:0] _RAND_41;
  reg [31:0] _RAND_42;
  reg [31:0] _RAND_43;
  reg [31:0] _RAND_44;
  reg [31:0] _RAND_45;
  reg [31:0] _RAND_46;
  reg [31:0] _RAND_47;
  reg [31:0] _RAND_48;
  reg [31:0] _RAND_49;
  reg [31:0] _RAND_50;
  reg [31:0] _RAND_51;
  reg [31:0] _RAND_52;
  reg [31:0] _RAND_53;
  reg [31:0] _RAND_54;
  reg [31:0] _RAND_55;
  reg [31:0] _RAND_56;
  reg [31:0] _RAND_57;
  reg [31:0] _RAND_58;
  reg [31:0] _RAND_59;
  reg [31:0] _RAND_60;
  reg [31:0] _RAND_61;
  reg [31:0] _RAND_62;
  reg [31:0] _RAND_63;
`endif // RANDOMIZE_REG_INIT
  reg [16:0] swdata_1_r_re; // @[Reg.scala 19:16]
  reg [16:0] swdata_1_r_im; // @[Reg.scala 19:16]
  reg [16:0] swdata_1_r_1_re; // @[Reg.scala 19:16]
  reg [16:0] swdata_1_r_1_im; // @[Reg.scala 19:16]
  reg [16:0] swdata_1_r_2_re; // @[Reg.scala 19:16]
  reg [16:0] swdata_1_r_2_im; // @[Reg.scala 19:16]
  reg [16:0] swdata_1_r_3_re; // @[Reg.scala 19:16]
  reg [16:0] swdata_1_r_3_im; // @[Reg.scala 19:16]
  reg [16:0] swdata_1_r_4_re; // @[Reg.scala 19:16]
  reg [16:0] swdata_1_r_4_im; // @[Reg.scala 19:16]
  reg [16:0] swdata_1_r_5_re; // @[Reg.scala 19:16]
  reg [16:0] swdata_1_r_5_im; // @[Reg.scala 19:16]
  reg [16:0] swdata_1_r_6_re; // @[Reg.scala 19:16]
  reg [16:0] swdata_1_r_6_im; // @[Reg.scala 19:16]
  reg [16:0] swdata_1_r_7_re; // @[Reg.scala 19:16]
  reg [16:0] swdata_1_r_7_im; // @[Reg.scala 19:16]
  reg [16:0] swdata_1_r_8_re; // @[Reg.scala 19:16]
  reg [16:0] swdata_1_r_8_im; // @[Reg.scala 19:16]
  reg [16:0] swdata_1_r_9_re; // @[Reg.scala 19:16]
  reg [16:0] swdata_1_r_9_im; // @[Reg.scala 19:16]
  reg [16:0] swdata_1_r_10_re; // @[Reg.scala 19:16]
  reg [16:0] swdata_1_r_10_im; // @[Reg.scala 19:16]
  reg [16:0] swdata_1_r_11_re; // @[Reg.scala 19:16]
  reg [16:0] swdata_1_r_11_im; // @[Reg.scala 19:16]
  reg [16:0] swdata_1_r_12_re; // @[Reg.scala 19:16]
  reg [16:0] swdata_1_r_12_im; // @[Reg.scala 19:16]
  reg [16:0] swdata_1_r_13_re; // @[Reg.scala 19:16]
  reg [16:0] swdata_1_r_13_im; // @[Reg.scala 19:16]
  reg [16:0] swdata_1_r_14_re; // @[Reg.scala 19:16]
  reg [16:0] swdata_1_r_14_im; // @[Reg.scala 19:16]
  reg [16:0] swdata_1_r_15_re; // @[Reg.scala 19:16]
  reg [16:0] swdata_1_r_15_im; // @[Reg.scala 19:16]
  reg [16:0] io_out_0_r_re; // @[Reg.scala 19:16]
  reg [16:0] io_out_0_r_im; // @[Reg.scala 19:16]
  reg [16:0] io_out_0_r_1_re; // @[Reg.scala 19:16]
  reg [16:0] io_out_0_r_1_im; // @[Reg.scala 19:16]
  reg [16:0] io_out_0_r_2_re; // @[Reg.scala 19:16]
  reg [16:0] io_out_0_r_2_im; // @[Reg.scala 19:16]
  reg [16:0] io_out_0_r_3_re; // @[Reg.scala 19:16]
  reg [16:0] io_out_0_r_3_im; // @[Reg.scala 19:16]
  reg [16:0] io_out_0_r_4_re; // @[Reg.scala 19:16]
  reg [16:0] io_out_0_r_4_im; // @[Reg.scala 19:16]
  reg [16:0] io_out_0_r_5_re; // @[Reg.scala 19:16]
  reg [16:0] io_out_0_r_5_im; // @[Reg.scala 19:16]
  reg [16:0] io_out_0_r_6_re; // @[Reg.scala 19:16]
  reg [16:0] io_out_0_r_6_im; // @[Reg.scala 19:16]
  reg [16:0] io_out_0_r_7_re; // @[Reg.scala 19:16]
  reg [16:0] io_out_0_r_7_im; // @[Reg.scala 19:16]
  reg [16:0] io_out_0_r_8_re; // @[Reg.scala 19:16]
  reg [16:0] io_out_0_r_8_im; // @[Reg.scala 19:16]
  reg [16:0] io_out_0_r_9_re; // @[Reg.scala 19:16]
  reg [16:0] io_out_0_r_9_im; // @[Reg.scala 19:16]
  reg [16:0] io_out_0_r_10_re; // @[Reg.scala 19:16]
  reg [16:0] io_out_0_r_10_im; // @[Reg.scala 19:16]
  reg [16:0] io_out_0_r_11_re; // @[Reg.scala 19:16]
  reg [16:0] io_out_0_r_11_im; // @[Reg.scala 19:16]
  reg [16:0] io_out_0_r_12_re; // @[Reg.scala 19:16]
  reg [16:0] io_out_0_r_12_im; // @[Reg.scala 19:16]
  reg [16:0] io_out_0_r_13_re; // @[Reg.scala 19:16]
  reg [16:0] io_out_0_r_13_im; // @[Reg.scala 19:16]
  reg [16:0] io_out_0_r_14_re; // @[Reg.scala 19:16]
  reg [16:0] io_out_0_r_14_im; // @[Reg.scala 19:16]
  reg [16:0] io_out_0_r_15_re; // @[Reg.scala 19:16]
  reg [16:0] io_out_0_r_15_im; // @[Reg.scala 19:16]
  assign io_out_0_re = io_out_0_r_15_re; // @[Modules.scala 306:38]
  assign io_out_0_im = io_out_0_r_15_im; // @[Modules.scala 306:38]
  assign io_out_1_re = io_sel ? io_in_0_re : swdata_1_r_15_re; // @[Modules.scala 306:{38,38}]
  assign io_out_1_im = io_sel ? io_in_0_im : swdata_1_r_15_im; // @[Modules.scala 306:{38,38}]
  always @(posedge clock) begin
    swdata_1_r_re <= io_in_1_re; // @[Reg.scala 19:16 20:{18,22}]
    swdata_1_r_im <= io_in_1_im; // @[Reg.scala 19:16 20:{18,22}]
    swdata_1_r_1_re <= swdata_1_r_re; // @[Reg.scala 19:16 20:{18,22}]
    swdata_1_r_1_im <= swdata_1_r_im; // @[Reg.scala 19:16 20:{18,22}]
    swdata_1_r_2_re <= swdata_1_r_1_re; // @[Reg.scala 19:16 20:{18,22}]
    swdata_1_r_2_im <= swdata_1_r_1_im; // @[Reg.scala 19:16 20:{18,22}]
    swdata_1_r_3_re <= swdata_1_r_2_re; // @[Reg.scala 19:16 20:{18,22}]
    swdata_1_r_3_im <= swdata_1_r_2_im; // @[Reg.scala 19:16 20:{18,22}]
    swdata_1_r_4_re <= swdata_1_r_3_re; // @[Reg.scala 19:16 20:{18,22}]
    swdata_1_r_4_im <= swdata_1_r_3_im; // @[Reg.scala 19:16 20:{18,22}]
    swdata_1_r_5_re <= swdata_1_r_4_re; // @[Reg.scala 19:16 20:{18,22}]
    swdata_1_r_5_im <= swdata_1_r_4_im; // @[Reg.scala 19:16 20:{18,22}]
    swdata_1_r_6_re <= swdata_1_r_5_re; // @[Reg.scala 19:16 20:{18,22}]
    swdata_1_r_6_im <= swdata_1_r_5_im; // @[Reg.scala 19:16 20:{18,22}]
    swdata_1_r_7_re <= swdata_1_r_6_re; // @[Reg.scala 19:16 20:{18,22}]
    swdata_1_r_7_im <= swdata_1_r_6_im; // @[Reg.scala 19:16 20:{18,22}]
    swdata_1_r_8_re <= swdata_1_r_7_re; // @[Reg.scala 19:16 20:{18,22}]
    swdata_1_r_8_im <= swdata_1_r_7_im; // @[Reg.scala 19:16 20:{18,22}]
    swdata_1_r_9_re <= swdata_1_r_8_re; // @[Reg.scala 19:16 20:{18,22}]
    swdata_1_r_9_im <= swdata_1_r_8_im; // @[Reg.scala 19:16 20:{18,22}]
    swdata_1_r_10_re <= swdata_1_r_9_re; // @[Reg.scala 19:16 20:{18,22}]
    swdata_1_r_10_im <= swdata_1_r_9_im; // @[Reg.scala 19:16 20:{18,22}]
    swdata_1_r_11_re <= swdata_1_r_10_re; // @[Reg.scala 19:16 20:{18,22}]
    swdata_1_r_11_im <= swdata_1_r_10_im; // @[Reg.scala 19:16 20:{18,22}]
    swdata_1_r_12_re <= swdata_1_r_11_re; // @[Reg.scala 19:16 20:{18,22}]
    swdata_1_r_12_im <= swdata_1_r_11_im; // @[Reg.scala 19:16 20:{18,22}]
    swdata_1_r_13_re <= swdata_1_r_12_re; // @[Reg.scala 19:16 20:{18,22}]
    swdata_1_r_13_im <= swdata_1_r_12_im; // @[Reg.scala 19:16 20:{18,22}]
    swdata_1_r_14_re <= swdata_1_r_13_re; // @[Reg.scala 19:16 20:{18,22}]
    swdata_1_r_14_im <= swdata_1_r_13_im; // @[Reg.scala 19:16 20:{18,22}]
    swdata_1_r_15_re <= swdata_1_r_14_re; // @[Reg.scala 19:16 20:{18,22}]
    swdata_1_r_15_im <= swdata_1_r_14_im; // @[Reg.scala 19:16 20:{18,22}]
    if (io_sel) begin // @[Reg.scala 20:22]
      io_out_0_r_re <= swdata_1_r_15_re; // @[Reg.scala 20:22]
    end else begin
      io_out_0_r_re <= io_in_0_re;
    end
    if (io_sel) begin // @[Reg.scala 20:22]
      io_out_0_r_im <= swdata_1_r_15_im; // @[Reg.scala 20:22]
    end else begin
      io_out_0_r_im <= io_in_0_im;
    end
    io_out_0_r_1_re <= io_out_0_r_re; // @[Reg.scala 19:16 20:{18,22}]
    io_out_0_r_1_im <= io_out_0_r_im; // @[Reg.scala 19:16 20:{18,22}]
    io_out_0_r_2_re <= io_out_0_r_1_re; // @[Reg.scala 19:16 20:{18,22}]
    io_out_0_r_2_im <= io_out_0_r_1_im; // @[Reg.scala 19:16 20:{18,22}]
    io_out_0_r_3_re <= io_out_0_r_2_re; // @[Reg.scala 19:16 20:{18,22}]
    io_out_0_r_3_im <= io_out_0_r_2_im; // @[Reg.scala 19:16 20:{18,22}]
    io_out_0_r_4_re <= io_out_0_r_3_re; // @[Reg.scala 19:16 20:{18,22}]
    io_out_0_r_4_im <= io_out_0_r_3_im; // @[Reg.scala 19:16 20:{18,22}]
    io_out_0_r_5_re <= io_out_0_r_4_re; // @[Reg.scala 19:16 20:{18,22}]
    io_out_0_r_5_im <= io_out_0_r_4_im; // @[Reg.scala 19:16 20:{18,22}]
    io_out_0_r_6_re <= io_out_0_r_5_re; // @[Reg.scala 19:16 20:{18,22}]
    io_out_0_r_6_im <= io_out_0_r_5_im; // @[Reg.scala 19:16 20:{18,22}]
    io_out_0_r_7_re <= io_out_0_r_6_re; // @[Reg.scala 19:16 20:{18,22}]
    io_out_0_r_7_im <= io_out_0_r_6_im; // @[Reg.scala 19:16 20:{18,22}]
    io_out_0_r_8_re <= io_out_0_r_7_re; // @[Reg.scala 19:16 20:{18,22}]
    io_out_0_r_8_im <= io_out_0_r_7_im; // @[Reg.scala 19:16 20:{18,22}]
    io_out_0_r_9_re <= io_out_0_r_8_re; // @[Reg.scala 19:16 20:{18,22}]
    io_out_0_r_9_im <= io_out_0_r_8_im; // @[Reg.scala 19:16 20:{18,22}]
    io_out_0_r_10_re <= io_out_0_r_9_re; // @[Reg.scala 19:16 20:{18,22}]
    io_out_0_r_10_im <= io_out_0_r_9_im; // @[Reg.scala 19:16 20:{18,22}]
    io_out_0_r_11_re <= io_out_0_r_10_re; // @[Reg.scala 19:16 20:{18,22}]
    io_out_0_r_11_im <= io_out_0_r_10_im; // @[Reg.scala 19:16 20:{18,22}]
    io_out_0_r_12_re <= io_out_0_r_11_re; // @[Reg.scala 19:16 20:{18,22}]
    io_out_0_r_12_im <= io_out_0_r_11_im; // @[Reg.scala 19:16 20:{18,22}]
    io_out_0_r_13_re <= io_out_0_r_12_re; // @[Reg.scala 19:16 20:{18,22}]
    io_out_0_r_13_im <= io_out_0_r_12_im; // @[Reg.scala 19:16 20:{18,22}]
    io_out_0_r_14_re <= io_out_0_r_13_re; // @[Reg.scala 19:16 20:{18,22}]
    io_out_0_r_14_im <= io_out_0_r_13_im; // @[Reg.scala 19:16 20:{18,22}]
    io_out_0_r_15_re <= io_out_0_r_14_re; // @[Reg.scala 19:16 20:{18,22}]
    io_out_0_r_15_im <= io_out_0_r_14_im; // @[Reg.scala 19:16 20:{18,22}]
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  swdata_1_r_re = _RAND_0[16:0];
  _RAND_1 = {1{`RANDOM}};
  swdata_1_r_im = _RAND_1[16:0];
  _RAND_2 = {1{`RANDOM}};
  swdata_1_r_1_re = _RAND_2[16:0];
  _RAND_3 = {1{`RANDOM}};
  swdata_1_r_1_im = _RAND_3[16:0];
  _RAND_4 = {1{`RANDOM}};
  swdata_1_r_2_re = _RAND_4[16:0];
  _RAND_5 = {1{`RANDOM}};
  swdata_1_r_2_im = _RAND_5[16:0];
  _RAND_6 = {1{`RANDOM}};
  swdata_1_r_3_re = _RAND_6[16:0];
  _RAND_7 = {1{`RANDOM}};
  swdata_1_r_3_im = _RAND_7[16:0];
  _RAND_8 = {1{`RANDOM}};
  swdata_1_r_4_re = _RAND_8[16:0];
  _RAND_9 = {1{`RANDOM}};
  swdata_1_r_4_im = _RAND_9[16:0];
  _RAND_10 = {1{`RANDOM}};
  swdata_1_r_5_re = _RAND_10[16:0];
  _RAND_11 = {1{`RANDOM}};
  swdata_1_r_5_im = _RAND_11[16:0];
  _RAND_12 = {1{`RANDOM}};
  swdata_1_r_6_re = _RAND_12[16:0];
  _RAND_13 = {1{`RANDOM}};
  swdata_1_r_6_im = _RAND_13[16:0];
  _RAND_14 = {1{`RANDOM}};
  swdata_1_r_7_re = _RAND_14[16:0];
  _RAND_15 = {1{`RANDOM}};
  swdata_1_r_7_im = _RAND_15[16:0];
  _RAND_16 = {1{`RANDOM}};
  swdata_1_r_8_re = _RAND_16[16:0];
  _RAND_17 = {1{`RANDOM}};
  swdata_1_r_8_im = _RAND_17[16:0];
  _RAND_18 = {1{`RANDOM}};
  swdata_1_r_9_re = _RAND_18[16:0];
  _RAND_19 = {1{`RANDOM}};
  swdata_1_r_9_im = _RAND_19[16:0];
  _RAND_20 = {1{`RANDOM}};
  swdata_1_r_10_re = _RAND_20[16:0];
  _RAND_21 = {1{`RANDOM}};
  swdata_1_r_10_im = _RAND_21[16:0];
  _RAND_22 = {1{`RANDOM}};
  swdata_1_r_11_re = _RAND_22[16:0];
  _RAND_23 = {1{`RANDOM}};
  swdata_1_r_11_im = _RAND_23[16:0];
  _RAND_24 = {1{`RANDOM}};
  swdata_1_r_12_re = _RAND_24[16:0];
  _RAND_25 = {1{`RANDOM}};
  swdata_1_r_12_im = _RAND_25[16:0];
  _RAND_26 = {1{`RANDOM}};
  swdata_1_r_13_re = _RAND_26[16:0];
  _RAND_27 = {1{`RANDOM}};
  swdata_1_r_13_im = _RAND_27[16:0];
  _RAND_28 = {1{`RANDOM}};
  swdata_1_r_14_re = _RAND_28[16:0];
  _RAND_29 = {1{`RANDOM}};
  swdata_1_r_14_im = _RAND_29[16:0];
  _RAND_30 = {1{`RANDOM}};
  swdata_1_r_15_re = _RAND_30[16:0];
  _RAND_31 = {1{`RANDOM}};
  swdata_1_r_15_im = _RAND_31[16:0];
  _RAND_32 = {1{`RANDOM}};
  io_out_0_r_re = _RAND_32[16:0];
  _RAND_33 = {1{`RANDOM}};
  io_out_0_r_im = _RAND_33[16:0];
  _RAND_34 = {1{`RANDOM}};
  io_out_0_r_1_re = _RAND_34[16:0];
  _RAND_35 = {1{`RANDOM}};
  io_out_0_r_1_im = _RAND_35[16:0];
  _RAND_36 = {1{`RANDOM}};
  io_out_0_r_2_re = _RAND_36[16:0];
  _RAND_37 = {1{`RANDOM}};
  io_out_0_r_2_im = _RAND_37[16:0];
  _RAND_38 = {1{`RANDOM}};
  io_out_0_r_3_re = _RAND_38[16:0];
  _RAND_39 = {1{`RANDOM}};
  io_out_0_r_3_im = _RAND_39[16:0];
  _RAND_40 = {1{`RANDOM}};
  io_out_0_r_4_re = _RAND_40[16:0];
  _RAND_41 = {1{`RANDOM}};
  io_out_0_r_4_im = _RAND_41[16:0];
  _RAND_42 = {1{`RANDOM}};
  io_out_0_r_5_re = _RAND_42[16:0];
  _RAND_43 = {1{`RANDOM}};
  io_out_0_r_5_im = _RAND_43[16:0];
  _RAND_44 = {1{`RANDOM}};
  io_out_0_r_6_re = _RAND_44[16:0];
  _RAND_45 = {1{`RANDOM}};
  io_out_0_r_6_im = _RAND_45[16:0];
  _RAND_46 = {1{`RANDOM}};
  io_out_0_r_7_re = _RAND_46[16:0];
  _RAND_47 = {1{`RANDOM}};
  io_out_0_r_7_im = _RAND_47[16:0];
  _RAND_48 = {1{`RANDOM}};
  io_out_0_r_8_re = _RAND_48[16:0];
  _RAND_49 = {1{`RANDOM}};
  io_out_0_r_8_im = _RAND_49[16:0];
  _RAND_50 = {1{`RANDOM}};
  io_out_0_r_9_re = _RAND_50[16:0];
  _RAND_51 = {1{`RANDOM}};
  io_out_0_r_9_im = _RAND_51[16:0];
  _RAND_52 = {1{`RANDOM}};
  io_out_0_r_10_re = _RAND_52[16:0];
  _RAND_53 = {1{`RANDOM}};
  io_out_0_r_10_im = _RAND_53[16:0];
  _RAND_54 = {1{`RANDOM}};
  io_out_0_r_11_re = _RAND_54[16:0];
  _RAND_55 = {1{`RANDOM}};
  io_out_0_r_11_im = _RAND_55[16:0];
  _RAND_56 = {1{`RANDOM}};
  io_out_0_r_12_re = _RAND_56[16:0];
  _RAND_57 = {1{`RANDOM}};
  io_out_0_r_12_im = _RAND_57[16:0];
  _RAND_58 = {1{`RANDOM}};
  io_out_0_r_13_re = _RAND_58[16:0];
  _RAND_59 = {1{`RANDOM}};
  io_out_0_r_13_im = _RAND_59[16:0];
  _RAND_60 = {1{`RANDOM}};
  io_out_0_r_14_re = _RAND_60[16:0];
  _RAND_61 = {1{`RANDOM}};
  io_out_0_r_14_im = _RAND_61[16:0];
  _RAND_62 = {1{`RANDOM}};
  io_out_0_r_15_re = _RAND_62[16:0];
  _RAND_63 = {1{`RANDOM}};
  io_out_0_r_15_im = _RAND_63[16:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module Switch_3(
  input         clock,
  input  [16:0] io_in_0_re,
  input  [16:0] io_in_0_im,
  input  [16:0] io_in_1_re,
  input  [16:0] io_in_1_im,
  output [16:0] io_out_0_re,
  output [16:0] io_out_0_im,
  output [16:0] io_out_1_re,
  output [16:0] io_out_1_im,
  input         io_sel
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_9;
  reg [31:0] _RAND_10;
  reg [31:0] _RAND_11;
  reg [31:0] _RAND_12;
  reg [31:0] _RAND_13;
  reg [31:0] _RAND_14;
  reg [31:0] _RAND_15;
  reg [31:0] _RAND_16;
  reg [31:0] _RAND_17;
  reg [31:0] _RAND_18;
  reg [31:0] _RAND_19;
  reg [31:0] _RAND_20;
  reg [31:0] _RAND_21;
  reg [31:0] _RAND_22;
  reg [31:0] _RAND_23;
  reg [31:0] _RAND_24;
  reg [31:0] _RAND_25;
  reg [31:0] _RAND_26;
  reg [31:0] _RAND_27;
  reg [31:0] _RAND_28;
  reg [31:0] _RAND_29;
  reg [31:0] _RAND_30;
  reg [31:0] _RAND_31;
`endif // RANDOMIZE_REG_INIT
  reg [16:0] swdata_1_r_re; // @[Reg.scala 19:16]
  reg [16:0] swdata_1_r_im; // @[Reg.scala 19:16]
  reg [16:0] swdata_1_r_1_re; // @[Reg.scala 19:16]
  reg [16:0] swdata_1_r_1_im; // @[Reg.scala 19:16]
  reg [16:0] swdata_1_r_2_re; // @[Reg.scala 19:16]
  reg [16:0] swdata_1_r_2_im; // @[Reg.scala 19:16]
  reg [16:0] swdata_1_r_3_re; // @[Reg.scala 19:16]
  reg [16:0] swdata_1_r_3_im; // @[Reg.scala 19:16]
  reg [16:0] swdata_1_r_4_re; // @[Reg.scala 19:16]
  reg [16:0] swdata_1_r_4_im; // @[Reg.scala 19:16]
  reg [16:0] swdata_1_r_5_re; // @[Reg.scala 19:16]
  reg [16:0] swdata_1_r_5_im; // @[Reg.scala 19:16]
  reg [16:0] swdata_1_r_6_re; // @[Reg.scala 19:16]
  reg [16:0] swdata_1_r_6_im; // @[Reg.scala 19:16]
  reg [16:0] swdata_1_r_7_re; // @[Reg.scala 19:16]
  reg [16:0] swdata_1_r_7_im; // @[Reg.scala 19:16]
  reg [16:0] io_out_0_r_re; // @[Reg.scala 19:16]
  reg [16:0] io_out_0_r_im; // @[Reg.scala 19:16]
  reg [16:0] io_out_0_r_1_re; // @[Reg.scala 19:16]
  reg [16:0] io_out_0_r_1_im; // @[Reg.scala 19:16]
  reg [16:0] io_out_0_r_2_re; // @[Reg.scala 19:16]
  reg [16:0] io_out_0_r_2_im; // @[Reg.scala 19:16]
  reg [16:0] io_out_0_r_3_re; // @[Reg.scala 19:16]
  reg [16:0] io_out_0_r_3_im; // @[Reg.scala 19:16]
  reg [16:0] io_out_0_r_4_re; // @[Reg.scala 19:16]
  reg [16:0] io_out_0_r_4_im; // @[Reg.scala 19:16]
  reg [16:0] io_out_0_r_5_re; // @[Reg.scala 19:16]
  reg [16:0] io_out_0_r_5_im; // @[Reg.scala 19:16]
  reg [16:0] io_out_0_r_6_re; // @[Reg.scala 19:16]
  reg [16:0] io_out_0_r_6_im; // @[Reg.scala 19:16]
  reg [16:0] io_out_0_r_7_re; // @[Reg.scala 19:16]
  reg [16:0] io_out_0_r_7_im; // @[Reg.scala 19:16]
  assign io_out_0_re = io_out_0_r_7_re; // @[Modules.scala 306:38]
  assign io_out_0_im = io_out_0_r_7_im; // @[Modules.scala 306:38]
  assign io_out_1_re = io_sel ? io_in_0_re : swdata_1_r_7_re; // @[Modules.scala 306:{38,38}]
  assign io_out_1_im = io_sel ? io_in_0_im : swdata_1_r_7_im; // @[Modules.scala 306:{38,38}]
  always @(posedge clock) begin
    swdata_1_r_re <= io_in_1_re; // @[Reg.scala 19:16 20:{18,22}]
    swdata_1_r_im <= io_in_1_im; // @[Reg.scala 19:16 20:{18,22}]
    swdata_1_r_1_re <= swdata_1_r_re; // @[Reg.scala 19:16 20:{18,22}]
    swdata_1_r_1_im <= swdata_1_r_im; // @[Reg.scala 19:16 20:{18,22}]
    swdata_1_r_2_re <= swdata_1_r_1_re; // @[Reg.scala 19:16 20:{18,22}]
    swdata_1_r_2_im <= swdata_1_r_1_im; // @[Reg.scala 19:16 20:{18,22}]
    swdata_1_r_3_re <= swdata_1_r_2_re; // @[Reg.scala 19:16 20:{18,22}]
    swdata_1_r_3_im <= swdata_1_r_2_im; // @[Reg.scala 19:16 20:{18,22}]
    swdata_1_r_4_re <= swdata_1_r_3_re; // @[Reg.scala 19:16 20:{18,22}]
    swdata_1_r_4_im <= swdata_1_r_3_im; // @[Reg.scala 19:16 20:{18,22}]
    swdata_1_r_5_re <= swdata_1_r_4_re; // @[Reg.scala 19:16 20:{18,22}]
    swdata_1_r_5_im <= swdata_1_r_4_im; // @[Reg.scala 19:16 20:{18,22}]
    swdata_1_r_6_re <= swdata_1_r_5_re; // @[Reg.scala 19:16 20:{18,22}]
    swdata_1_r_6_im <= swdata_1_r_5_im; // @[Reg.scala 19:16 20:{18,22}]
    swdata_1_r_7_re <= swdata_1_r_6_re; // @[Reg.scala 19:16 20:{18,22}]
    swdata_1_r_7_im <= swdata_1_r_6_im; // @[Reg.scala 19:16 20:{18,22}]
    if (io_sel) begin // @[Reg.scala 20:22]
      io_out_0_r_re <= swdata_1_r_7_re; // @[Reg.scala 20:22]
    end else begin
      io_out_0_r_re <= io_in_0_re;
    end
    if (io_sel) begin // @[Reg.scala 20:22]
      io_out_0_r_im <= swdata_1_r_7_im; // @[Reg.scala 20:22]
    end else begin
      io_out_0_r_im <= io_in_0_im;
    end
    io_out_0_r_1_re <= io_out_0_r_re; // @[Reg.scala 19:16 20:{18,22}]
    io_out_0_r_1_im <= io_out_0_r_im; // @[Reg.scala 19:16 20:{18,22}]
    io_out_0_r_2_re <= io_out_0_r_1_re; // @[Reg.scala 19:16 20:{18,22}]
    io_out_0_r_2_im <= io_out_0_r_1_im; // @[Reg.scala 19:16 20:{18,22}]
    io_out_0_r_3_re <= io_out_0_r_2_re; // @[Reg.scala 19:16 20:{18,22}]
    io_out_0_r_3_im <= io_out_0_r_2_im; // @[Reg.scala 19:16 20:{18,22}]
    io_out_0_r_4_re <= io_out_0_r_3_re; // @[Reg.scala 19:16 20:{18,22}]
    io_out_0_r_4_im <= io_out_0_r_3_im; // @[Reg.scala 19:16 20:{18,22}]
    io_out_0_r_5_re <= io_out_0_r_4_re; // @[Reg.scala 19:16 20:{18,22}]
    io_out_0_r_5_im <= io_out_0_r_4_im; // @[Reg.scala 19:16 20:{18,22}]
    io_out_0_r_6_re <= io_out_0_r_5_re; // @[Reg.scala 19:16 20:{18,22}]
    io_out_0_r_6_im <= io_out_0_r_5_im; // @[Reg.scala 19:16 20:{18,22}]
    io_out_0_r_7_re <= io_out_0_r_6_re; // @[Reg.scala 19:16 20:{18,22}]
    io_out_0_r_7_im <= io_out_0_r_6_im; // @[Reg.scala 19:16 20:{18,22}]
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  swdata_1_r_re = _RAND_0[16:0];
  _RAND_1 = {1{`RANDOM}};
  swdata_1_r_im = _RAND_1[16:0];
  _RAND_2 = {1{`RANDOM}};
  swdata_1_r_1_re = _RAND_2[16:0];
  _RAND_3 = {1{`RANDOM}};
  swdata_1_r_1_im = _RAND_3[16:0];
  _RAND_4 = {1{`RANDOM}};
  swdata_1_r_2_re = _RAND_4[16:0];
  _RAND_5 = {1{`RANDOM}};
  swdata_1_r_2_im = _RAND_5[16:0];
  _RAND_6 = {1{`RANDOM}};
  swdata_1_r_3_re = _RAND_6[16:0];
  _RAND_7 = {1{`RANDOM}};
  swdata_1_r_3_im = _RAND_7[16:0];
  _RAND_8 = {1{`RANDOM}};
  swdata_1_r_4_re = _RAND_8[16:0];
  _RAND_9 = {1{`RANDOM}};
  swdata_1_r_4_im = _RAND_9[16:0];
  _RAND_10 = {1{`RANDOM}};
  swdata_1_r_5_re = _RAND_10[16:0];
  _RAND_11 = {1{`RANDOM}};
  swdata_1_r_5_im = _RAND_11[16:0];
  _RAND_12 = {1{`RANDOM}};
  swdata_1_r_6_re = _RAND_12[16:0];
  _RAND_13 = {1{`RANDOM}};
  swdata_1_r_6_im = _RAND_13[16:0];
  _RAND_14 = {1{`RANDOM}};
  swdata_1_r_7_re = _RAND_14[16:0];
  _RAND_15 = {1{`RANDOM}};
  swdata_1_r_7_im = _RAND_15[16:0];
  _RAND_16 = {1{`RANDOM}};
  io_out_0_r_re = _RAND_16[16:0];
  _RAND_17 = {1{`RANDOM}};
  io_out_0_r_im = _RAND_17[16:0];
  _RAND_18 = {1{`RANDOM}};
  io_out_0_r_1_re = _RAND_18[16:0];
  _RAND_19 = {1{`RANDOM}};
  io_out_0_r_1_im = _RAND_19[16:0];
  _RAND_20 = {1{`RANDOM}};
  io_out_0_r_2_re = _RAND_20[16:0];
  _RAND_21 = {1{`RANDOM}};
  io_out_0_r_2_im = _RAND_21[16:0];
  _RAND_22 = {1{`RANDOM}};
  io_out_0_r_3_re = _RAND_22[16:0];
  _RAND_23 = {1{`RANDOM}};
  io_out_0_r_3_im = _RAND_23[16:0];
  _RAND_24 = {1{`RANDOM}};
  io_out_0_r_4_re = _RAND_24[16:0];
  _RAND_25 = {1{`RANDOM}};
  io_out_0_r_4_im = _RAND_25[16:0];
  _RAND_26 = {1{`RANDOM}};
  io_out_0_r_5_re = _RAND_26[16:0];
  _RAND_27 = {1{`RANDOM}};
  io_out_0_r_5_im = _RAND_27[16:0];
  _RAND_28 = {1{`RANDOM}};
  io_out_0_r_6_re = _RAND_28[16:0];
  _RAND_29 = {1{`RANDOM}};
  io_out_0_r_6_im = _RAND_29[16:0];
  _RAND_30 = {1{`RANDOM}};
  io_out_0_r_7_re = _RAND_30[16:0];
  _RAND_31 = {1{`RANDOM}};
  io_out_0_r_7_im = _RAND_31[16:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module Switch_4(
  input         clock,
  input  [16:0] io_in_0_re,
  input  [16:0] io_in_0_im,
  input  [16:0] io_in_1_re,
  input  [16:0] io_in_1_im,
  output [16:0] io_out_0_re,
  output [16:0] io_out_0_im,
  output [16:0] io_out_1_re,
  output [16:0] io_out_1_im,
  input         io_sel
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_9;
  reg [31:0] _RAND_10;
  reg [31:0] _RAND_11;
  reg [31:0] _RAND_12;
  reg [31:0] _RAND_13;
  reg [31:0] _RAND_14;
  reg [31:0] _RAND_15;
`endif // RANDOMIZE_REG_INIT
  reg [16:0] swdata_1_r_re; // @[Reg.scala 19:16]
  reg [16:0] swdata_1_r_im; // @[Reg.scala 19:16]
  reg [16:0] swdata_1_r_1_re; // @[Reg.scala 19:16]
  reg [16:0] swdata_1_r_1_im; // @[Reg.scala 19:16]
  reg [16:0] swdata_1_r_2_re; // @[Reg.scala 19:16]
  reg [16:0] swdata_1_r_2_im; // @[Reg.scala 19:16]
  reg [16:0] swdata_1_r_3_re; // @[Reg.scala 19:16]
  reg [16:0] swdata_1_r_3_im; // @[Reg.scala 19:16]
  reg [16:0] io_out_0_r_re; // @[Reg.scala 19:16]
  reg [16:0] io_out_0_r_im; // @[Reg.scala 19:16]
  reg [16:0] io_out_0_r_1_re; // @[Reg.scala 19:16]
  reg [16:0] io_out_0_r_1_im; // @[Reg.scala 19:16]
  reg [16:0] io_out_0_r_2_re; // @[Reg.scala 19:16]
  reg [16:0] io_out_0_r_2_im; // @[Reg.scala 19:16]
  reg [16:0] io_out_0_r_3_re; // @[Reg.scala 19:16]
  reg [16:0] io_out_0_r_3_im; // @[Reg.scala 19:16]
  assign io_out_0_re = io_out_0_r_3_re; // @[Modules.scala 306:38]
  assign io_out_0_im = io_out_0_r_3_im; // @[Modules.scala 306:38]
  assign io_out_1_re = io_sel ? io_in_0_re : swdata_1_r_3_re; // @[Modules.scala 306:{38,38}]
  assign io_out_1_im = io_sel ? io_in_0_im : swdata_1_r_3_im; // @[Modules.scala 306:{38,38}]
  always @(posedge clock) begin
    swdata_1_r_re <= io_in_1_re; // @[Reg.scala 19:16 20:{18,22}]
    swdata_1_r_im <= io_in_1_im; // @[Reg.scala 19:16 20:{18,22}]
    swdata_1_r_1_re <= swdata_1_r_re; // @[Reg.scala 19:16 20:{18,22}]
    swdata_1_r_1_im <= swdata_1_r_im; // @[Reg.scala 19:16 20:{18,22}]
    swdata_1_r_2_re <= swdata_1_r_1_re; // @[Reg.scala 19:16 20:{18,22}]
    swdata_1_r_2_im <= swdata_1_r_1_im; // @[Reg.scala 19:16 20:{18,22}]
    swdata_1_r_3_re <= swdata_1_r_2_re; // @[Reg.scala 19:16 20:{18,22}]
    swdata_1_r_3_im <= swdata_1_r_2_im; // @[Reg.scala 19:16 20:{18,22}]
    if (io_sel) begin // @[Reg.scala 20:22]
      io_out_0_r_re <= swdata_1_r_3_re; // @[Reg.scala 20:22]
    end else begin
      io_out_0_r_re <= io_in_0_re;
    end
    if (io_sel) begin // @[Reg.scala 20:22]
      io_out_0_r_im <= swdata_1_r_3_im; // @[Reg.scala 20:22]
    end else begin
      io_out_0_r_im <= io_in_0_im;
    end
    io_out_0_r_1_re <= io_out_0_r_re; // @[Reg.scala 19:16 20:{18,22}]
    io_out_0_r_1_im <= io_out_0_r_im; // @[Reg.scala 19:16 20:{18,22}]
    io_out_0_r_2_re <= io_out_0_r_1_re; // @[Reg.scala 19:16 20:{18,22}]
    io_out_0_r_2_im <= io_out_0_r_1_im; // @[Reg.scala 19:16 20:{18,22}]
    io_out_0_r_3_re <= io_out_0_r_2_re; // @[Reg.scala 19:16 20:{18,22}]
    io_out_0_r_3_im <= io_out_0_r_2_im; // @[Reg.scala 19:16 20:{18,22}]
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  swdata_1_r_re = _RAND_0[16:0];
  _RAND_1 = {1{`RANDOM}};
  swdata_1_r_im = _RAND_1[16:0];
  _RAND_2 = {1{`RANDOM}};
  swdata_1_r_1_re = _RAND_2[16:0];
  _RAND_3 = {1{`RANDOM}};
  swdata_1_r_1_im = _RAND_3[16:0];
  _RAND_4 = {1{`RANDOM}};
  swdata_1_r_2_re = _RAND_4[16:0];
  _RAND_5 = {1{`RANDOM}};
  swdata_1_r_2_im = _RAND_5[16:0];
  _RAND_6 = {1{`RANDOM}};
  swdata_1_r_3_re = _RAND_6[16:0];
  _RAND_7 = {1{`RANDOM}};
  swdata_1_r_3_im = _RAND_7[16:0];
  _RAND_8 = {1{`RANDOM}};
  io_out_0_r_re = _RAND_8[16:0];
  _RAND_9 = {1{`RANDOM}};
  io_out_0_r_im = _RAND_9[16:0];
  _RAND_10 = {1{`RANDOM}};
  io_out_0_r_1_re = _RAND_10[16:0];
  _RAND_11 = {1{`RANDOM}};
  io_out_0_r_1_im = _RAND_11[16:0];
  _RAND_12 = {1{`RANDOM}};
  io_out_0_r_2_re = _RAND_12[16:0];
  _RAND_13 = {1{`RANDOM}};
  io_out_0_r_2_im = _RAND_13[16:0];
  _RAND_14 = {1{`RANDOM}};
  io_out_0_r_3_re = _RAND_14[16:0];
  _RAND_15 = {1{`RANDOM}};
  io_out_0_r_3_im = _RAND_15[16:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module Switch_5(
  input         clock,
  input  [16:0] io_in_0_re,
  input  [16:0] io_in_0_im,
  input  [16:0] io_in_1_re,
  input  [16:0] io_in_1_im,
  output [16:0] io_out_0_re,
  output [16:0] io_out_0_im,
  output [16:0] io_out_1_re,
  output [16:0] io_out_1_im,
  input         io_sel
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
`endif // RANDOMIZE_REG_INIT
  reg [16:0] swdata_1_r_re; // @[Reg.scala 19:16]
  reg [16:0] swdata_1_r_im; // @[Reg.scala 19:16]
  reg [16:0] swdata_1_r_1_re; // @[Reg.scala 19:16]
  reg [16:0] swdata_1_r_1_im; // @[Reg.scala 19:16]
  reg [16:0] io_out_0_r_re; // @[Reg.scala 19:16]
  reg [16:0] io_out_0_r_im; // @[Reg.scala 19:16]
  reg [16:0] io_out_0_r_1_re; // @[Reg.scala 19:16]
  reg [16:0] io_out_0_r_1_im; // @[Reg.scala 19:16]
  assign io_out_0_re = io_out_0_r_1_re; // @[Modules.scala 306:38]
  assign io_out_0_im = io_out_0_r_1_im; // @[Modules.scala 306:38]
  assign io_out_1_re = io_sel ? io_in_0_re : swdata_1_r_1_re; // @[Modules.scala 306:{38,38}]
  assign io_out_1_im = io_sel ? io_in_0_im : swdata_1_r_1_im; // @[Modules.scala 306:{38,38}]
  always @(posedge clock) begin
    swdata_1_r_re <= io_in_1_re; // @[Reg.scala 19:16 20:{18,22}]
    swdata_1_r_im <= io_in_1_im; // @[Reg.scala 19:16 20:{18,22}]
    swdata_1_r_1_re <= swdata_1_r_re; // @[Reg.scala 19:16 20:{18,22}]
    swdata_1_r_1_im <= swdata_1_r_im; // @[Reg.scala 19:16 20:{18,22}]
    if (io_sel) begin // @[Reg.scala 20:22]
      io_out_0_r_re <= swdata_1_r_1_re; // @[Reg.scala 20:22]
    end else begin
      io_out_0_r_re <= io_in_0_re;
    end
    if (io_sel) begin // @[Reg.scala 20:22]
      io_out_0_r_im <= swdata_1_r_1_im; // @[Reg.scala 20:22]
    end else begin
      io_out_0_r_im <= io_in_0_im;
    end
    io_out_0_r_1_re <= io_out_0_r_re; // @[Reg.scala 19:16 20:{18,22}]
    io_out_0_r_1_im <= io_out_0_r_im; // @[Reg.scala 19:16 20:{18,22}]
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  swdata_1_r_re = _RAND_0[16:0];
  _RAND_1 = {1{`RANDOM}};
  swdata_1_r_im = _RAND_1[16:0];
  _RAND_2 = {1{`RANDOM}};
  swdata_1_r_1_re = _RAND_2[16:0];
  _RAND_3 = {1{`RANDOM}};
  swdata_1_r_1_im = _RAND_3[16:0];
  _RAND_4 = {1{`RANDOM}};
  io_out_0_r_re = _RAND_4[16:0];
  _RAND_5 = {1{`RANDOM}};
  io_out_0_r_im = _RAND_5[16:0];
  _RAND_6 = {1{`RANDOM}};
  io_out_0_r_1_re = _RAND_6[16:0];
  _RAND_7 = {1{`RANDOM}};
  io_out_0_r_1_im = _RAND_7[16:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module Switch_6(
  input         clock,
  input  [16:0] io_in_0_re,
  input  [16:0] io_in_0_im,
  input  [16:0] io_in_1_re,
  input  [16:0] io_in_1_im,
  output [16:0] io_out_0_re,
  output [16:0] io_out_0_im,
  output [16:0] io_out_1_re,
  output [16:0] io_out_1_im,
  input         io_sel
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
`endif // RANDOMIZE_REG_INIT
  reg [16:0] swdata_1_r_re; // @[Reg.scala 19:16]
  reg [16:0] swdata_1_r_im; // @[Reg.scala 19:16]
  reg [16:0] io_out_0_r_re; // @[Reg.scala 19:16]
  reg [16:0] io_out_0_r_im; // @[Reg.scala 19:16]
  assign io_out_0_re = io_out_0_r_re; // @[Modules.scala 306:38]
  assign io_out_0_im = io_out_0_r_im; // @[Modules.scala 306:38]
  assign io_out_1_re = io_sel ? io_in_0_re : swdata_1_r_re; // @[Modules.scala 306:{38,38}]
  assign io_out_1_im = io_sel ? io_in_0_im : swdata_1_r_im; // @[Modules.scala 306:{38,38}]
  always @(posedge clock) begin
    swdata_1_r_re <= io_in_1_re; // @[Reg.scala 19:16 20:{18,22}]
    swdata_1_r_im <= io_in_1_im; // @[Reg.scala 19:16 20:{18,22}]
    if (io_sel) begin // @[Reg.scala 20:22]
      io_out_0_r_re <= swdata_1_r_re; // @[Reg.scala 20:22]
    end else begin
      io_out_0_r_re <= io_in_0_re;
    end
    if (io_sel) begin // @[Reg.scala 20:22]
      io_out_0_r_im <= swdata_1_r_im; // @[Reg.scala 20:22]
    end else begin
      io_out_0_r_im <= io_in_0_im;
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  swdata_1_r_re = _RAND_0[16:0];
  _RAND_1 = {1{`RANDOM}};
  swdata_1_r_im = _RAND_1[16:0];
  _RAND_2 = {1{`RANDOM}};
  io_out_0_r_re = _RAND_2[16:0];
  _RAND_3 = {1{`RANDOM}};
  io_out_0_r_im = _RAND_3[16:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module ComplexRecode(
  input  [15:0] io_in_re,
  input  [15:0] io_in_im,
  output [16:0] io_out_re,
  output [16:0] io_out_im
);
  wire  io_out_re_rawIn_sign = io_in_re[15]; // @[rawFloatFromFN.scala 46:22]
  wire [4:0] io_out_re_rawIn_expIn = io_in_re[14:10]; // @[rawFloatFromFN.scala 47:23]
  wire [9:0] io_out_re_rawIn_fractIn = io_in_re[9:0]; // @[rawFloatFromFN.scala 48:25]
  wire  io_out_re_rawIn_isZeroExpIn = io_out_re_rawIn_expIn == 5'h0; // @[rawFloatFromFN.scala 50:34]
  wire  io_out_re_rawIn_isZeroFractIn = io_out_re_rawIn_fractIn == 10'h0; // @[rawFloatFromFN.scala 51:38]
  wire [3:0] _io_out_re_rawIn_normDist_T_10 = io_out_re_rawIn_fractIn[1] ? 4'h8 : 4'h9; // @[Mux.scala 47:70]
  wire [3:0] _io_out_re_rawIn_normDist_T_11 = io_out_re_rawIn_fractIn[2] ? 4'h7 : _io_out_re_rawIn_normDist_T_10; // @[Mux.scala 47:70]
  wire [3:0] _io_out_re_rawIn_normDist_T_12 = io_out_re_rawIn_fractIn[3] ? 4'h6 : _io_out_re_rawIn_normDist_T_11; // @[Mux.scala 47:70]
  wire [3:0] _io_out_re_rawIn_normDist_T_13 = io_out_re_rawIn_fractIn[4] ? 4'h5 : _io_out_re_rawIn_normDist_T_12; // @[Mux.scala 47:70]
  wire [3:0] _io_out_re_rawIn_normDist_T_14 = io_out_re_rawIn_fractIn[5] ? 4'h4 : _io_out_re_rawIn_normDist_T_13; // @[Mux.scala 47:70]
  wire [3:0] _io_out_re_rawIn_normDist_T_15 = io_out_re_rawIn_fractIn[6] ? 4'h3 : _io_out_re_rawIn_normDist_T_14; // @[Mux.scala 47:70]
  wire [3:0] _io_out_re_rawIn_normDist_T_16 = io_out_re_rawIn_fractIn[7] ? 4'h2 : _io_out_re_rawIn_normDist_T_15; // @[Mux.scala 47:70]
  wire [3:0] _io_out_re_rawIn_normDist_T_17 = io_out_re_rawIn_fractIn[8] ? 4'h1 : _io_out_re_rawIn_normDist_T_16; // @[Mux.scala 47:70]
  wire [3:0] io_out_re_rawIn_normDist = io_out_re_rawIn_fractIn[9] ? 4'h0 : _io_out_re_rawIn_normDist_T_17; // @[Mux.scala 47:70]
  wire [24:0] _GEN_8 = {{15'd0}, io_out_re_rawIn_fractIn}; // @[rawFloatFromFN.scala 54:36]
  wire [24:0] _io_out_re_rawIn_subnormFract_T = _GEN_8 << io_out_re_rawIn_normDist; // @[rawFloatFromFN.scala 54:36]
  wire [9:0] io_out_re_rawIn_subnormFract = {_io_out_re_rawIn_subnormFract_T[8:0], 1'h0}; // @[rawFloatFromFN.scala 54:64]
  wire [5:0] _GEN_0 = {{2'd0}, io_out_re_rawIn_normDist}; // @[rawFloatFromFN.scala 57:26]
  wire [5:0] _io_out_re_rawIn_adjustedExp_T = _GEN_0 ^ 6'h3f; // @[rawFloatFromFN.scala 57:26]
  wire [5:0] _io_out_re_rawIn_adjustedExp_T_1 = io_out_re_rawIn_isZeroExpIn ? _io_out_re_rawIn_adjustedExp_T : {{1'd0},
    io_out_re_rawIn_expIn}; // @[rawFloatFromFN.scala 56:16]
  wire [1:0] _io_out_re_rawIn_adjustedExp_T_2 = io_out_re_rawIn_isZeroExpIn ? 2'h2 : 2'h1; // @[rawFloatFromFN.scala 60:27]
  wire [4:0] _GEN_1 = {{3'd0}, _io_out_re_rawIn_adjustedExp_T_2}; // @[rawFloatFromFN.scala 60:22]
  wire [4:0] _io_out_re_rawIn_adjustedExp_T_3 = 5'h10 | _GEN_1; // @[rawFloatFromFN.scala 60:22]
  wire [5:0] _GEN_2 = {{1'd0}, _io_out_re_rawIn_adjustedExp_T_3}; // @[rawFloatFromFN.scala 59:15]
  wire [5:0] io_out_re_rawIn_adjustedExp = _io_out_re_rawIn_adjustedExp_T_1 + _GEN_2; // @[rawFloatFromFN.scala 59:15]
  wire  io_out_re_rawIn_isZero = io_out_re_rawIn_isZeroExpIn & io_out_re_rawIn_isZeroFractIn; // @[rawFloatFromFN.scala 62:34]
  wire  io_out_re_rawIn_isSpecial = io_out_re_rawIn_adjustedExp[5:4] == 2'h3; // @[rawFloatFromFN.scala 63:62]
  wire  io_out_re_rawIn__isNaN = io_out_re_rawIn_isSpecial & ~io_out_re_rawIn_isZeroFractIn; // @[rawFloatFromFN.scala 66:33]
  wire [6:0] io_out_re_rawIn__sExp = {1'b0,$signed(io_out_re_rawIn_adjustedExp)}; // @[rawFloatFromFN.scala 70:48]
  wire  _io_out_re_rawIn_out_sig_T = ~io_out_re_rawIn_isZero; // @[rawFloatFromFN.scala 72:29]
  wire [9:0] _io_out_re_rawIn_out_sig_T_1 = io_out_re_rawIn_isZeroExpIn ? io_out_re_rawIn_subnormFract :
    io_out_re_rawIn_fractIn; // @[rawFloatFromFN.scala 72:42]
  wire [11:0] io_out_re_rawIn__sig = {1'h0,_io_out_re_rawIn_out_sig_T,_io_out_re_rawIn_out_sig_T_1}; // @[Cat.scala 33:92]
  wire [2:0] _io_out_re_T_1 = io_out_re_rawIn_isZero ? 3'h0 : io_out_re_rawIn__sExp[5:3]; // @[recFNFromFN.scala 48:16]
  wire [2:0] _GEN_3 = {{2'd0}, io_out_re_rawIn__isNaN}; // @[recFNFromFN.scala 48:79]
  wire [2:0] _io_out_re_T_3 = _io_out_re_T_1 | _GEN_3; // @[recFNFromFN.scala 48:79]
  wire [12:0] io_out_re_lo = {io_out_re_rawIn__sExp[2:0],io_out_re_rawIn__sig[9:0]}; // @[Cat.scala 33:92]
  wire [3:0] io_out_re_hi = {io_out_re_rawIn_sign,_io_out_re_T_3}; // @[Cat.scala 33:92]
  wire  io_out_im_rawIn_sign = io_in_im[15]; // @[rawFloatFromFN.scala 46:22]
  wire [4:0] io_out_im_rawIn_expIn = io_in_im[14:10]; // @[rawFloatFromFN.scala 47:23]
  wire [9:0] io_out_im_rawIn_fractIn = io_in_im[9:0]; // @[rawFloatFromFN.scala 48:25]
  wire  io_out_im_rawIn_isZeroExpIn = io_out_im_rawIn_expIn == 5'h0; // @[rawFloatFromFN.scala 50:34]
  wire  io_out_im_rawIn_isZeroFractIn = io_out_im_rawIn_fractIn == 10'h0; // @[rawFloatFromFN.scala 51:38]
  wire [3:0] _io_out_im_rawIn_normDist_T_10 = io_out_im_rawIn_fractIn[1] ? 4'h8 : 4'h9; // @[Mux.scala 47:70]
  wire [3:0] _io_out_im_rawIn_normDist_T_11 = io_out_im_rawIn_fractIn[2] ? 4'h7 : _io_out_im_rawIn_normDist_T_10; // @[Mux.scala 47:70]
  wire [3:0] _io_out_im_rawIn_normDist_T_12 = io_out_im_rawIn_fractIn[3] ? 4'h6 : _io_out_im_rawIn_normDist_T_11; // @[Mux.scala 47:70]
  wire [3:0] _io_out_im_rawIn_normDist_T_13 = io_out_im_rawIn_fractIn[4] ? 4'h5 : _io_out_im_rawIn_normDist_T_12; // @[Mux.scala 47:70]
  wire [3:0] _io_out_im_rawIn_normDist_T_14 = io_out_im_rawIn_fractIn[5] ? 4'h4 : _io_out_im_rawIn_normDist_T_13; // @[Mux.scala 47:70]
  wire [3:0] _io_out_im_rawIn_normDist_T_15 = io_out_im_rawIn_fractIn[6] ? 4'h3 : _io_out_im_rawIn_normDist_T_14; // @[Mux.scala 47:70]
  wire [3:0] _io_out_im_rawIn_normDist_T_16 = io_out_im_rawIn_fractIn[7] ? 4'h2 : _io_out_im_rawIn_normDist_T_15; // @[Mux.scala 47:70]
  wire [3:0] _io_out_im_rawIn_normDist_T_17 = io_out_im_rawIn_fractIn[8] ? 4'h1 : _io_out_im_rawIn_normDist_T_16; // @[Mux.scala 47:70]
  wire [3:0] io_out_im_rawIn_normDist = io_out_im_rawIn_fractIn[9] ? 4'h0 : _io_out_im_rawIn_normDist_T_17; // @[Mux.scala 47:70]
  wire [24:0] _GEN_9 = {{15'd0}, io_out_im_rawIn_fractIn}; // @[rawFloatFromFN.scala 54:36]
  wire [24:0] _io_out_im_rawIn_subnormFract_T = _GEN_9 << io_out_im_rawIn_normDist; // @[rawFloatFromFN.scala 54:36]
  wire [9:0] io_out_im_rawIn_subnormFract = {_io_out_im_rawIn_subnormFract_T[8:0], 1'h0}; // @[rawFloatFromFN.scala 54:64]
  wire [5:0] _GEN_4 = {{2'd0}, io_out_im_rawIn_normDist}; // @[rawFloatFromFN.scala 57:26]
  wire [5:0] _io_out_im_rawIn_adjustedExp_T = _GEN_4 ^ 6'h3f; // @[rawFloatFromFN.scala 57:26]
  wire [5:0] _io_out_im_rawIn_adjustedExp_T_1 = io_out_im_rawIn_isZeroExpIn ? _io_out_im_rawIn_adjustedExp_T : {{1'd0},
    io_out_im_rawIn_expIn}; // @[rawFloatFromFN.scala 56:16]
  wire [1:0] _io_out_im_rawIn_adjustedExp_T_2 = io_out_im_rawIn_isZeroExpIn ? 2'h2 : 2'h1; // @[rawFloatFromFN.scala 60:27]
  wire [4:0] _GEN_5 = {{3'd0}, _io_out_im_rawIn_adjustedExp_T_2}; // @[rawFloatFromFN.scala 60:22]
  wire [4:0] _io_out_im_rawIn_adjustedExp_T_3 = 5'h10 | _GEN_5; // @[rawFloatFromFN.scala 60:22]
  wire [5:0] _GEN_6 = {{1'd0}, _io_out_im_rawIn_adjustedExp_T_3}; // @[rawFloatFromFN.scala 59:15]
  wire [5:0] io_out_im_rawIn_adjustedExp = _io_out_im_rawIn_adjustedExp_T_1 + _GEN_6; // @[rawFloatFromFN.scala 59:15]
  wire  io_out_im_rawIn_isZero = io_out_im_rawIn_isZeroExpIn & io_out_im_rawIn_isZeroFractIn; // @[rawFloatFromFN.scala 62:34]
  wire  io_out_im_rawIn_isSpecial = io_out_im_rawIn_adjustedExp[5:4] == 2'h3; // @[rawFloatFromFN.scala 63:62]
  wire  io_out_im_rawIn__isNaN = io_out_im_rawIn_isSpecial & ~io_out_im_rawIn_isZeroFractIn; // @[rawFloatFromFN.scala 66:33]
  wire [6:0] io_out_im_rawIn__sExp = {1'b0,$signed(io_out_im_rawIn_adjustedExp)}; // @[rawFloatFromFN.scala 70:48]
  wire  _io_out_im_rawIn_out_sig_T = ~io_out_im_rawIn_isZero; // @[rawFloatFromFN.scala 72:29]
  wire [9:0] _io_out_im_rawIn_out_sig_T_1 = io_out_im_rawIn_isZeroExpIn ? io_out_im_rawIn_subnormFract :
    io_out_im_rawIn_fractIn; // @[rawFloatFromFN.scala 72:42]
  wire [11:0] io_out_im_rawIn__sig = {1'h0,_io_out_im_rawIn_out_sig_T,_io_out_im_rawIn_out_sig_T_1}; // @[Cat.scala 33:92]
  wire [2:0] _io_out_im_T_1 = io_out_im_rawIn_isZero ? 3'h0 : io_out_im_rawIn__sExp[5:3]; // @[recFNFromFN.scala 48:16]
  wire [2:0] _GEN_7 = {{2'd0}, io_out_im_rawIn__isNaN}; // @[recFNFromFN.scala 48:79]
  wire [2:0] _io_out_im_T_3 = _io_out_im_T_1 | _GEN_7; // @[recFNFromFN.scala 48:79]
  wire [12:0] io_out_im_lo = {io_out_im_rawIn__sExp[2:0],io_out_im_rawIn__sig[9:0]}; // @[Cat.scala 33:92]
  wire [3:0] io_out_im_hi = {io_out_im_rawIn_sign,_io_out_im_T_3}; // @[Cat.scala 33:92]
  assign io_out_re = {io_out_re_hi,io_out_re_lo}; // @[Cat.scala 33:92]
  assign io_out_im = {io_out_im_hi,io_out_im_lo}; // @[Cat.scala 33:92]
endmodule
module ComplexDecode(
  input  [16:0] io_in_re,
  input  [16:0] io_in_im,
  output [15:0] io_out_re,
  output [15:0] io_out_im
);
  wire [5:0] io_out_re_rawIn_exp = io_in_re[15:10]; // @[rawFloatFromRecFN.scala 50:21]
  wire  io_out_re_rawIn_isZero = io_out_re_rawIn_exp[5:3] == 3'h0; // @[rawFloatFromRecFN.scala 51:54]
  wire  io_out_re_rawIn_isSpecial = io_out_re_rawIn_exp[5:4] == 2'h3; // @[rawFloatFromRecFN.scala 52:54]
  wire  io_out_re_rawIn__isNaN = io_out_re_rawIn_isSpecial & io_out_re_rawIn_exp[3]; // @[rawFloatFromRecFN.scala 55:33]
  wire  io_out_re_rawIn__isInf = io_out_re_rawIn_isSpecial & ~io_out_re_rawIn_exp[3]; // @[rawFloatFromRecFN.scala 56:33]
  wire  io_out_re_rawIn__sign = io_in_re[16]; // @[rawFloatFromRecFN.scala 58:25]
  wire [6:0] io_out_re_rawIn__sExp = {1'b0,$signed(io_out_re_rawIn_exp)}; // @[rawFloatFromRecFN.scala 59:27]
  wire  _io_out_re_rawIn_out_sig_T = ~io_out_re_rawIn_isZero; // @[rawFloatFromRecFN.scala 60:39]
  wire [11:0] io_out_re_rawIn__sig = {1'h0,_io_out_re_rawIn_out_sig_T,io_in_re[9:0]}; // @[Cat.scala 33:92]
  wire  io_out_re_isSubnormal = $signed(io_out_re_rawIn__sExp) < 7'sh12; // @[fNFromRecFN.scala 50:39]
  wire [3:0] io_out_re_denormShiftDist = 4'h1 - io_out_re_rawIn__sExp[3:0]; // @[fNFromRecFN.scala 51:39]
  wire [10:0] _io_out_re_denormFract_T_1 = io_out_re_rawIn__sig[11:1] >> io_out_re_denormShiftDist; // @[fNFromRecFN.scala 52:42]
  wire [9:0] io_out_re_denormFract = _io_out_re_denormFract_T_1[9:0]; // @[fNFromRecFN.scala 52:60]
  wire [4:0] _io_out_re_expOut_T_2 = io_out_re_rawIn__sExp[4:0] - 5'h11; // @[fNFromRecFN.scala 57:45]
  wire [4:0] _io_out_re_expOut_T_3 = io_out_re_isSubnormal ? 5'h0 : _io_out_re_expOut_T_2; // @[fNFromRecFN.scala 55:16]
  wire  _io_out_re_expOut_T_4 = io_out_re_rawIn__isNaN | io_out_re_rawIn__isInf; // @[fNFromRecFN.scala 59:44]
  wire [4:0] _io_out_re_expOut_T_6 = _io_out_re_expOut_T_4 ? 5'h1f : 5'h0; // @[Bitwise.scala 77:12]
  wire [4:0] io_out_re_expOut = _io_out_re_expOut_T_3 | _io_out_re_expOut_T_6; // @[fNFromRecFN.scala 59:15]
  wire [9:0] _io_out_re_fractOut_T_1 = io_out_re_rawIn__isInf ? 10'h0 : io_out_re_rawIn__sig[9:0]; // @[fNFromRecFN.scala 63:20]
  wire [9:0] io_out_re_fractOut = io_out_re_isSubnormal ? io_out_re_denormFract : _io_out_re_fractOut_T_1; // @[fNFromRecFN.scala 61:16]
  wire [5:0] io_out_re_hi = {io_out_re_rawIn__sign,io_out_re_expOut}; // @[Cat.scala 33:92]
  wire [5:0] io_out_im_rawIn_exp = io_in_im[15:10]; // @[rawFloatFromRecFN.scala 50:21]
  wire  io_out_im_rawIn_isZero = io_out_im_rawIn_exp[5:3] == 3'h0; // @[rawFloatFromRecFN.scala 51:54]
  wire  io_out_im_rawIn_isSpecial = io_out_im_rawIn_exp[5:4] == 2'h3; // @[rawFloatFromRecFN.scala 52:54]
  wire  io_out_im_rawIn__isNaN = io_out_im_rawIn_isSpecial & io_out_im_rawIn_exp[3]; // @[rawFloatFromRecFN.scala 55:33]
  wire  io_out_im_rawIn__isInf = io_out_im_rawIn_isSpecial & ~io_out_im_rawIn_exp[3]; // @[rawFloatFromRecFN.scala 56:33]
  wire  io_out_im_rawIn__sign = io_in_im[16]; // @[rawFloatFromRecFN.scala 58:25]
  wire [6:0] io_out_im_rawIn__sExp = {1'b0,$signed(io_out_im_rawIn_exp)}; // @[rawFloatFromRecFN.scala 59:27]
  wire  _io_out_im_rawIn_out_sig_T = ~io_out_im_rawIn_isZero; // @[rawFloatFromRecFN.scala 60:39]
  wire [11:0] io_out_im_rawIn__sig = {1'h0,_io_out_im_rawIn_out_sig_T,io_in_im[9:0]}; // @[Cat.scala 33:92]
  wire  io_out_im_isSubnormal = $signed(io_out_im_rawIn__sExp) < 7'sh12; // @[fNFromRecFN.scala 50:39]
  wire [3:0] io_out_im_denormShiftDist = 4'h1 - io_out_im_rawIn__sExp[3:0]; // @[fNFromRecFN.scala 51:39]
  wire [10:0] _io_out_im_denormFract_T_1 = io_out_im_rawIn__sig[11:1] >> io_out_im_denormShiftDist; // @[fNFromRecFN.scala 52:42]
  wire [9:0] io_out_im_denormFract = _io_out_im_denormFract_T_1[9:0]; // @[fNFromRecFN.scala 52:60]
  wire [4:0] _io_out_im_expOut_T_2 = io_out_im_rawIn__sExp[4:0] - 5'h11; // @[fNFromRecFN.scala 57:45]
  wire [4:0] _io_out_im_expOut_T_3 = io_out_im_isSubnormal ? 5'h0 : _io_out_im_expOut_T_2; // @[fNFromRecFN.scala 55:16]
  wire  _io_out_im_expOut_T_4 = io_out_im_rawIn__isNaN | io_out_im_rawIn__isInf; // @[fNFromRecFN.scala 59:44]
  wire [4:0] _io_out_im_expOut_T_6 = _io_out_im_expOut_T_4 ? 5'h1f : 5'h0; // @[Bitwise.scala 77:12]
  wire [4:0] io_out_im_expOut = _io_out_im_expOut_T_3 | _io_out_im_expOut_T_6; // @[fNFromRecFN.scala 59:15]
  wire [9:0] _io_out_im_fractOut_T_1 = io_out_im_rawIn__isInf ? 10'h0 : io_out_im_rawIn__sig[9:0]; // @[fNFromRecFN.scala 63:20]
  wire [9:0] io_out_im_fractOut = io_out_im_isSubnormal ? io_out_im_denormFract : _io_out_im_fractOut_T_1; // @[fNFromRecFN.scala 61:16]
  wire [5:0] io_out_im_hi = {io_out_im_rawIn__sign,io_out_im_expOut}; // @[Cat.scala 33:92]
  assign io_out_re = {io_out_re_hi,io_out_re_fractOut}; // @[Cat.scala 33:92]
  assign io_out_im = {io_out_im_hi,io_out_im_fractOut}; // @[Cat.scala 33:92]
endmodule
module FFT(
  input         clock,
  input         reset,
  input  [15:0] io_dIn_0_re,
  input  [15:0] io_dIn_0_im,
  input  [15:0] io_dIn_1_re,
  input  [15:0] io_dIn_1_im,
  output [15:0] io_dOut_0_re,
  output [15:0] io_dOut_0_im,
  output [15:0] io_dOut_1_re,
  output [15:0] io_dOut_1_im,
  input         io_din_valid,
  output        io_dout_valid,
  output        io_busy
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
`endif // RANDOMIZE_REG_INIT
  wire [16:0] inst_io_in_0_re; // @[Modules.scala 287:22]
  wire [16:0] inst_io_in_0_im; // @[Modules.scala 287:22]
  wire [16:0] inst_io_in_1_re; // @[Modules.scala 287:22]
  wire [16:0] inst_io_in_1_im; // @[Modules.scala 287:22]
  wire [16:0] inst_io_out_0_re; // @[Modules.scala 287:22]
  wire [16:0] inst_io_out_0_im; // @[Modules.scala 287:22]
  wire [16:0] inst_io_out_1_re; // @[Modules.scala 287:22]
  wire [16:0] inst_io_out_1_im; // @[Modules.scala 287:22]
  wire [16:0] inst_io_wn_0_re; // @[Modules.scala 287:22]
  wire [16:0] inst_io_wn_0_im; // @[Modules.scala 287:22]
  wire [16:0] inst_1_io_in_0_re; // @[Modules.scala 287:22]
  wire [16:0] inst_1_io_in_0_im; // @[Modules.scala 287:22]
  wire [16:0] inst_1_io_in_1_re; // @[Modules.scala 287:22]
  wire [16:0] inst_1_io_in_1_im; // @[Modules.scala 287:22]
  wire [16:0] inst_1_io_out_0_re; // @[Modules.scala 287:22]
  wire [16:0] inst_1_io_out_0_im; // @[Modules.scala 287:22]
  wire [16:0] inst_1_io_out_1_re; // @[Modules.scala 287:22]
  wire [16:0] inst_1_io_out_1_im; // @[Modules.scala 287:22]
  wire [16:0] inst_1_io_wn_0_re; // @[Modules.scala 287:22]
  wire [16:0] inst_1_io_wn_0_im; // @[Modules.scala 287:22]
  wire [16:0] inst_2_io_in_0_re; // @[Modules.scala 287:22]
  wire [16:0] inst_2_io_in_0_im; // @[Modules.scala 287:22]
  wire [16:0] inst_2_io_in_1_re; // @[Modules.scala 287:22]
  wire [16:0] inst_2_io_in_1_im; // @[Modules.scala 287:22]
  wire [16:0] inst_2_io_out_0_re; // @[Modules.scala 287:22]
  wire [16:0] inst_2_io_out_0_im; // @[Modules.scala 287:22]
  wire [16:0] inst_2_io_out_1_re; // @[Modules.scala 287:22]
  wire [16:0] inst_2_io_out_1_im; // @[Modules.scala 287:22]
  wire [16:0] inst_2_io_wn_0_re; // @[Modules.scala 287:22]
  wire [16:0] inst_2_io_wn_0_im; // @[Modules.scala 287:22]
  wire [16:0] inst_3_io_in_0_re; // @[Modules.scala 287:22]
  wire [16:0] inst_3_io_in_0_im; // @[Modules.scala 287:22]
  wire [16:0] inst_3_io_in_1_re; // @[Modules.scala 287:22]
  wire [16:0] inst_3_io_in_1_im; // @[Modules.scala 287:22]
  wire [16:0] inst_3_io_out_0_re; // @[Modules.scala 287:22]
  wire [16:0] inst_3_io_out_0_im; // @[Modules.scala 287:22]
  wire [16:0] inst_3_io_out_1_re; // @[Modules.scala 287:22]
  wire [16:0] inst_3_io_out_1_im; // @[Modules.scala 287:22]
  wire [16:0] inst_3_io_wn_0_re; // @[Modules.scala 287:22]
  wire [16:0] inst_3_io_wn_0_im; // @[Modules.scala 287:22]
  wire [16:0] inst_4_io_in_0_re; // @[Modules.scala 287:22]
  wire [16:0] inst_4_io_in_0_im; // @[Modules.scala 287:22]
  wire [16:0] inst_4_io_in_1_re; // @[Modules.scala 287:22]
  wire [16:0] inst_4_io_in_1_im; // @[Modules.scala 287:22]
  wire [16:0] inst_4_io_out_0_re; // @[Modules.scala 287:22]
  wire [16:0] inst_4_io_out_0_im; // @[Modules.scala 287:22]
  wire [16:0] inst_4_io_out_1_re; // @[Modules.scala 287:22]
  wire [16:0] inst_4_io_out_1_im; // @[Modules.scala 287:22]
  wire [16:0] inst_4_io_wn_0_re; // @[Modules.scala 287:22]
  wire [16:0] inst_4_io_wn_0_im; // @[Modules.scala 287:22]
  wire [16:0] inst_5_io_in_0_re; // @[Modules.scala 287:22]
  wire [16:0] inst_5_io_in_0_im; // @[Modules.scala 287:22]
  wire [16:0] inst_5_io_in_1_re; // @[Modules.scala 287:22]
  wire [16:0] inst_5_io_in_1_im; // @[Modules.scala 287:22]
  wire [16:0] inst_5_io_out_0_re; // @[Modules.scala 287:22]
  wire [16:0] inst_5_io_out_0_im; // @[Modules.scala 287:22]
  wire [16:0] inst_5_io_out_1_re; // @[Modules.scala 287:22]
  wire [16:0] inst_5_io_out_1_im; // @[Modules.scala 287:22]
  wire [16:0] inst_5_io_wn_0_re; // @[Modules.scala 287:22]
  wire [16:0] inst_5_io_wn_0_im; // @[Modules.scala 287:22]
  wire [16:0] inst_6_io_in_0_re; // @[Modules.scala 287:22]
  wire [16:0] inst_6_io_in_0_im; // @[Modules.scala 287:22]
  wire [16:0] inst_6_io_in_1_re; // @[Modules.scala 287:22]
  wire [16:0] inst_6_io_in_1_im; // @[Modules.scala 287:22]
  wire [16:0] inst_6_io_out_0_re; // @[Modules.scala 287:22]
  wire [16:0] inst_6_io_out_0_im; // @[Modules.scala 287:22]
  wire [16:0] inst_6_io_out_1_re; // @[Modules.scala 287:22]
  wire [16:0] inst_6_io_out_1_im; // @[Modules.scala 287:22]
  wire [16:0] inst_6_io_wn_0_re; // @[Modules.scala 287:22]
  wire [16:0] inst_6_io_wn_0_im; // @[Modules.scala 287:22]
  wire [16:0] dataotemp_inst_io_in_0_re; // @[Modules.scala 213:22]
  wire [16:0] dataotemp_inst_io_in_0_im; // @[Modules.scala 213:22]
  wire [16:0] dataotemp_inst_io_in_1_re; // @[Modules.scala 213:22]
  wire [16:0] dataotemp_inst_io_in_1_im; // @[Modules.scala 213:22]
  wire [16:0] dataotemp_inst_io_out_0_re; // @[Modules.scala 213:22]
  wire [16:0] dataotemp_inst_io_out_0_im; // @[Modules.scala 213:22]
  wire [16:0] dataotemp_inst_io_out_1_re; // @[Modules.scala 213:22]
  wire [16:0] dataotemp_inst_io_out_1_im; // @[Modules.scala 213:22]
  wire  inst_7_clock; // @[Modules.scala 311:22]
  wire [16:0] inst_7_io_in_0_re; // @[Modules.scala 311:22]
  wire [16:0] inst_7_io_in_0_im; // @[Modules.scala 311:22]
  wire [16:0] inst_7_io_in_1_re; // @[Modules.scala 311:22]
  wire [16:0] inst_7_io_in_1_im; // @[Modules.scala 311:22]
  wire [16:0] inst_7_io_out_0_re; // @[Modules.scala 311:22]
  wire [16:0] inst_7_io_out_0_im; // @[Modules.scala 311:22]
  wire [16:0] inst_7_io_out_1_re; // @[Modules.scala 311:22]
  wire [16:0] inst_7_io_out_1_im; // @[Modules.scala 311:22]
  wire  inst_7_io_sel; // @[Modules.scala 311:22]
  wire  inst_8_clock; // @[Modules.scala 311:22]
  wire [16:0] inst_8_io_in_0_re; // @[Modules.scala 311:22]
  wire [16:0] inst_8_io_in_0_im; // @[Modules.scala 311:22]
  wire [16:0] inst_8_io_in_1_re; // @[Modules.scala 311:22]
  wire [16:0] inst_8_io_in_1_im; // @[Modules.scala 311:22]
  wire [16:0] inst_8_io_out_0_re; // @[Modules.scala 311:22]
  wire [16:0] inst_8_io_out_0_im; // @[Modules.scala 311:22]
  wire [16:0] inst_8_io_out_1_re; // @[Modules.scala 311:22]
  wire [16:0] inst_8_io_out_1_im; // @[Modules.scala 311:22]
  wire  inst_8_io_sel; // @[Modules.scala 311:22]
  wire  inst_9_clock; // @[Modules.scala 311:22]
  wire [16:0] inst_9_io_in_0_re; // @[Modules.scala 311:22]
  wire [16:0] inst_9_io_in_0_im; // @[Modules.scala 311:22]
  wire [16:0] inst_9_io_in_1_re; // @[Modules.scala 311:22]
  wire [16:0] inst_9_io_in_1_im; // @[Modules.scala 311:22]
  wire [16:0] inst_9_io_out_0_re; // @[Modules.scala 311:22]
  wire [16:0] inst_9_io_out_0_im; // @[Modules.scala 311:22]
  wire [16:0] inst_9_io_out_1_re; // @[Modules.scala 311:22]
  wire [16:0] inst_9_io_out_1_im; // @[Modules.scala 311:22]
  wire  inst_9_io_sel; // @[Modules.scala 311:22]
  wire  inst_10_clock; // @[Modules.scala 311:22]
  wire [16:0] inst_10_io_in_0_re; // @[Modules.scala 311:22]
  wire [16:0] inst_10_io_in_0_im; // @[Modules.scala 311:22]
  wire [16:0] inst_10_io_in_1_re; // @[Modules.scala 311:22]
  wire [16:0] inst_10_io_in_1_im; // @[Modules.scala 311:22]
  wire [16:0] inst_10_io_out_0_re; // @[Modules.scala 311:22]
  wire [16:0] inst_10_io_out_0_im; // @[Modules.scala 311:22]
  wire [16:0] inst_10_io_out_1_re; // @[Modules.scala 311:22]
  wire [16:0] inst_10_io_out_1_im; // @[Modules.scala 311:22]
  wire  inst_10_io_sel; // @[Modules.scala 311:22]
  wire  inst_11_clock; // @[Modules.scala 311:22]
  wire [16:0] inst_11_io_in_0_re; // @[Modules.scala 311:22]
  wire [16:0] inst_11_io_in_0_im; // @[Modules.scala 311:22]
  wire [16:0] inst_11_io_in_1_re; // @[Modules.scala 311:22]
  wire [16:0] inst_11_io_in_1_im; // @[Modules.scala 311:22]
  wire [16:0] inst_11_io_out_0_re; // @[Modules.scala 311:22]
  wire [16:0] inst_11_io_out_0_im; // @[Modules.scala 311:22]
  wire [16:0] inst_11_io_out_1_re; // @[Modules.scala 311:22]
  wire [16:0] inst_11_io_out_1_im; // @[Modules.scala 311:22]
  wire  inst_11_io_sel; // @[Modules.scala 311:22]
  wire  inst_12_clock; // @[Modules.scala 311:22]
  wire [16:0] inst_12_io_in_0_re; // @[Modules.scala 311:22]
  wire [16:0] inst_12_io_in_0_im; // @[Modules.scala 311:22]
  wire [16:0] inst_12_io_in_1_re; // @[Modules.scala 311:22]
  wire [16:0] inst_12_io_in_1_im; // @[Modules.scala 311:22]
  wire [16:0] inst_12_io_out_0_re; // @[Modules.scala 311:22]
  wire [16:0] inst_12_io_out_0_im; // @[Modules.scala 311:22]
  wire [16:0] inst_12_io_out_1_re; // @[Modules.scala 311:22]
  wire [16:0] inst_12_io_out_1_im; // @[Modules.scala 311:22]
  wire  inst_12_io_sel; // @[Modules.scala 311:22]
  wire  inst_13_clock; // @[Modules.scala 311:22]
  wire [16:0] inst_13_io_in_0_re; // @[Modules.scala 311:22]
  wire [16:0] inst_13_io_in_0_im; // @[Modules.scala 311:22]
  wire [16:0] inst_13_io_in_1_re; // @[Modules.scala 311:22]
  wire [16:0] inst_13_io_in_1_im; // @[Modules.scala 311:22]
  wire [16:0] inst_13_io_out_0_re; // @[Modules.scala 311:22]
  wire [16:0] inst_13_io_out_0_im; // @[Modules.scala 311:22]
  wire [16:0] inst_13_io_out_1_re; // @[Modules.scala 311:22]
  wire [16:0] inst_13_io_out_1_im; // @[Modules.scala 311:22]
  wire  inst_13_io_sel; // @[Modules.scala 311:22]
  wire [15:0] inst_14_io_in_re; // @[Modules.scala 40:22]
  wire [15:0] inst_14_io_in_im; // @[Modules.scala 40:22]
  wire [16:0] inst_14_io_out_re; // @[Modules.scala 40:22]
  wire [16:0] inst_14_io_out_im; // @[Modules.scala 40:22]
  wire [15:0] inst_15_io_in_re; // @[Modules.scala 40:22]
  wire [15:0] inst_15_io_in_im; // @[Modules.scala 40:22]
  wire [16:0] inst_15_io_out_re; // @[Modules.scala 40:22]
  wire [16:0] inst_15_io_out_im; // @[Modules.scala 40:22]
  wire [16:0] inst_16_io_in_re; // @[Modules.scala 56:22]
  wire [16:0] inst_16_io_in_im; // @[Modules.scala 56:22]
  wire [15:0] inst_16_io_out_re; // @[Modules.scala 56:22]
  wire [15:0] inst_16_io_out_im; // @[Modules.scala 56:22]
  wire [16:0] inst_17_io_in_re; // @[Modules.scala 56:22]
  wire [16:0] inst_17_io_in_im; // @[Modules.scala 56:22]
  wire [15:0] inst_17_io_out_re; // @[Modules.scala 56:22]
  wire [15:0] inst_17_io_out_im; // @[Modules.scala 56:22]
  reg [8:0] cnt_0; // @[FFT.scala 110:46]
  wire  busy = cnt_0 != 9'h0; // @[FFT.scala 114:21]
  wire [8:0] _cnt_0_T_2 = cnt_0 + 9'h1; // @[FFT.scala 116:87]
  wire [6:0] wnCtrl = cnt_0[6:0]; // @[FFT.scala 131:23]
  wire [7:0] _wnList_T = {{1'd0}, wnCtrl}; // @[FFT.scala 135:96]
  wire [6:0] wnList_res_re_rawIn__sExp = {1'b0,$signed(6'h20)}; // @[rawFloatFromFN.scala 70:48]
  wire [16:0] _wnList_res_re_T_7 = {1'h0,wnList_res_re_rawIn__sExp[5:3],wnList_res_re_rawIn__sExp[2:0],10'h0}; // @[Cat.scala 33:92]
  wire [6:0] wnList_res_re_rawIn_1_sExp = {1'b0,$signed(6'h1f)}; // @[rawFloatFromFN.scala 70:48]
  wire [16:0] _wnList_res_re_T_15 = {1'h0,wnList_res_re_rawIn_1_sExp[5:3],wnList_res_re_rawIn_1_sExp[2:0],10'h3ff}; // @[Cat.scala 33:92]
  wire [16:0] _wnList_res_re_T_23 = {1'h0,wnList_res_re_rawIn_1_sExp[5:3],wnList_res_re_rawIn_1_sExp[2:0],10'h3fd}; // @[Cat.scala 33:92]
  wire [16:0] _wnList_res_re_T_31 = {1'h0,wnList_res_re_rawIn_1_sExp[5:3],wnList_res_re_rawIn_1_sExp[2:0],10'h3fa}; // @[Cat.scala 33:92]
  wire [16:0] _wnList_res_re_T_39 = {1'h0,wnList_res_re_rawIn_1_sExp[5:3],wnList_res_re_rawIn_1_sExp[2:0],10'h3f6}; // @[Cat.scala 33:92]
  wire [16:0] _wnList_res_re_T_47 = {1'h0,wnList_res_re_rawIn_1_sExp[5:3],wnList_res_re_rawIn_1_sExp[2:0],10'h3f0}; // @[Cat.scala 33:92]
  wire [16:0] _wnList_res_re_T_55 = {1'h0,wnList_res_re_rawIn_1_sExp[5:3],wnList_res_re_rawIn_1_sExp[2:0],10'h3e9}; // @[Cat.scala 33:92]
  wire [16:0] _wnList_res_re_T_63 = {1'h0,wnList_res_re_rawIn_1_sExp[5:3],wnList_res_re_rawIn_1_sExp[2:0],10'h3e1}; // @[Cat.scala 33:92]
  wire [16:0] _wnList_res_re_T_71 = {1'h0,wnList_res_re_rawIn_1_sExp[5:3],wnList_res_re_rawIn_1_sExp[2:0],10'h3d8}; // @[Cat.scala 33:92]
  wire [16:0] _wnList_res_re_T_79 = {1'h0,wnList_res_re_rawIn_1_sExp[5:3],wnList_res_re_rawIn_1_sExp[2:0],10'h3ce}; // @[Cat.scala 33:92]
  wire [16:0] _wnList_res_re_T_87 = {1'h0,wnList_res_re_rawIn_1_sExp[5:3],wnList_res_re_rawIn_1_sExp[2:0],10'h3c2}; // @[Cat.scala 33:92]
  wire [16:0] _wnList_res_re_T_95 = {1'h0,wnList_res_re_rawIn_1_sExp[5:3],wnList_res_re_rawIn_1_sExp[2:0],10'h3b5}; // @[Cat.scala 33:92]
  wire [16:0] _wnList_res_re_T_103 = {1'h0,wnList_res_re_rawIn_1_sExp[5:3],wnList_res_re_rawIn_1_sExp[2:0],10'h3a7}; // @[Cat.scala 33:92]
  wire [16:0] _wnList_res_re_T_111 = {1'h0,wnList_res_re_rawIn_1_sExp[5:3],wnList_res_re_rawIn_1_sExp[2:0],10'h398}; // @[Cat.scala 33:92]
  wire [16:0] _wnList_res_re_T_119 = {1'h0,wnList_res_re_rawIn_1_sExp[5:3],wnList_res_re_rawIn_1_sExp[2:0],10'h388}; // @[Cat.scala 33:92]
  wire [16:0] _wnList_res_re_T_127 = {1'h0,wnList_res_re_rawIn_1_sExp[5:3],wnList_res_re_rawIn_1_sExp[2:0],10'h376}; // @[Cat.scala 33:92]
  wire [16:0] _wnList_res_re_T_135 = {1'h0,wnList_res_re_rawIn_1_sExp[5:3],wnList_res_re_rawIn_1_sExp[2:0],10'h364}; // @[Cat.scala 33:92]
  wire [16:0] _wnList_res_re_T_143 = {1'h0,wnList_res_re_rawIn_1_sExp[5:3],wnList_res_re_rawIn_1_sExp[2:0],10'h350}; // @[Cat.scala 33:92]
  wire [16:0] _wnList_res_re_T_151 = {1'h0,wnList_res_re_rawIn_1_sExp[5:3],wnList_res_re_rawIn_1_sExp[2:0],10'h33b}; // @[Cat.scala 33:92]
  wire [16:0] _wnList_res_re_T_159 = {1'h0,wnList_res_re_rawIn_1_sExp[5:3],wnList_res_re_rawIn_1_sExp[2:0],10'h325}; // @[Cat.scala 33:92]
  wire [16:0] _wnList_res_re_T_167 = {1'h0,wnList_res_re_rawIn_1_sExp[5:3],wnList_res_re_rawIn_1_sExp[2:0],10'h30e}; // @[Cat.scala 33:92]
  wire [16:0] _wnList_res_re_T_175 = {1'h0,wnList_res_re_rawIn_1_sExp[5:3],wnList_res_re_rawIn_1_sExp[2:0],10'h2f5}; // @[Cat.scala 33:92]
  wire [16:0] _wnList_res_re_T_183 = {1'h0,wnList_res_re_rawIn_1_sExp[5:3],wnList_res_re_rawIn_1_sExp[2:0],10'h2dc}; // @[Cat.scala 33:92]
  wire [16:0] _wnList_res_re_T_191 = {1'h0,wnList_res_re_rawIn_1_sExp[5:3],wnList_res_re_rawIn_1_sExp[2:0],10'h2c2}; // @[Cat.scala 33:92]
  wire [16:0] _wnList_res_re_T_199 = {1'h0,wnList_res_re_rawIn_1_sExp[5:3],wnList_res_re_rawIn_1_sExp[2:0],10'h2a6}; // @[Cat.scala 33:92]
  wire [16:0] _wnList_res_re_T_207 = {1'h0,wnList_res_re_rawIn_1_sExp[5:3],wnList_res_re_rawIn_1_sExp[2:0],10'h28a}; // @[Cat.scala 33:92]
  wire [16:0] _wnList_res_re_T_215 = {1'h0,wnList_res_re_rawIn_1_sExp[5:3],wnList_res_re_rawIn_1_sExp[2:0],10'h26c}; // @[Cat.scala 33:92]
  wire [16:0] _wnList_res_re_T_223 = {1'h0,wnList_res_re_rawIn_1_sExp[5:3],wnList_res_re_rawIn_1_sExp[2:0],10'h24e}; // @[Cat.scala 33:92]
  wire [16:0] _wnList_res_re_T_231 = {1'h0,wnList_res_re_rawIn_1_sExp[5:3],wnList_res_re_rawIn_1_sExp[2:0],10'h22f}; // @[Cat.scala 33:92]
  wire [16:0] _wnList_res_re_T_239 = {1'h0,wnList_res_re_rawIn_1_sExp[5:3],wnList_res_re_rawIn_1_sExp[2:0],10'h20e}; // @[Cat.scala 33:92]
  wire [16:0] _wnList_res_re_T_247 = {1'h0,wnList_res_re_rawIn_1_sExp[5:3],wnList_res_re_rawIn_1_sExp[2:0],10'h1ed}; // @[Cat.scala 33:92]
  wire [16:0] _wnList_res_re_T_255 = {1'h0,wnList_res_re_rawIn_1_sExp[5:3],wnList_res_re_rawIn_1_sExp[2:0],10'h1cb}; // @[Cat.scala 33:92]
  wire [16:0] _wnList_res_re_T_263 = {1'h0,wnList_res_re_rawIn_1_sExp[5:3],wnList_res_re_rawIn_1_sExp[2:0],10'h1a8}; // @[Cat.scala 33:92]
  wire [16:0] _wnList_res_re_T_271 = {1'h0,wnList_res_re_rawIn_1_sExp[5:3],wnList_res_re_rawIn_1_sExp[2:0],10'h184}; // @[Cat.scala 33:92]
  wire [16:0] _wnList_res_re_T_279 = {1'h0,wnList_res_re_rawIn_1_sExp[5:3],wnList_res_re_rawIn_1_sExp[2:0],10'h15f}; // @[Cat.scala 33:92]
  wire [16:0] _wnList_res_re_T_287 = {1'h0,wnList_res_re_rawIn_1_sExp[5:3],wnList_res_re_rawIn_1_sExp[2:0],10'h139}; // @[Cat.scala 33:92]
  wire [16:0] _wnList_res_re_T_295 = {1'h0,wnList_res_re_rawIn_1_sExp[5:3],wnList_res_re_rawIn_1_sExp[2:0],10'h113}; // @[Cat.scala 33:92]
  wire [16:0] _wnList_res_re_T_303 = {1'h0,wnList_res_re_rawIn_1_sExp[5:3],wnList_res_re_rawIn_1_sExp[2:0],10'heb}; // @[Cat.scala 33:92]
  wire [16:0] _wnList_res_re_T_311 = {1'h0,wnList_res_re_rawIn_1_sExp[5:3],wnList_res_re_rawIn_1_sExp[2:0],10'hc3}; // @[Cat.scala 33:92]
  wire [16:0] _wnList_res_re_T_319 = {1'h0,wnList_res_re_rawIn_1_sExp[5:3],wnList_res_re_rawIn_1_sExp[2:0],10'h9b}; // @[Cat.scala 33:92]
  wire [16:0] _wnList_res_re_T_327 = {1'h0,wnList_res_re_rawIn_1_sExp[5:3],wnList_res_re_rawIn_1_sExp[2:0],10'h71}; // @[Cat.scala 33:92]
  wire [16:0] _wnList_res_re_T_335 = {1'h0,wnList_res_re_rawIn_1_sExp[5:3],wnList_res_re_rawIn_1_sExp[2:0],10'h47}; // @[Cat.scala 33:92]
  wire [16:0] _wnList_res_re_T_343 = {1'h0,wnList_res_re_rawIn_1_sExp[5:3],wnList_res_re_rawIn_1_sExp[2:0],10'h1c}; // @[Cat.scala 33:92]
  wire [6:0] wnList_res_re_rawIn_43_sExp = {1'b0,$signed(6'h1e)}; // @[rawFloatFromFN.scala 70:48]
  wire [16:0] _wnList_res_re_T_351 = {1'h0,wnList_res_re_rawIn_43_sExp[5:3],wnList_res_re_rawIn_43_sExp[2:0],10'h3e2}; // @[Cat.scala 33:92]
  wire [16:0] _wnList_res_re_T_359 = {1'h0,wnList_res_re_rawIn_43_sExp[5:3],wnList_res_re_rawIn_43_sExp[2:0],10'h38a}; // @[Cat.scala 33:92]
  wire [16:0] _wnList_res_re_T_367 = {1'h0,wnList_res_re_rawIn_43_sExp[5:3],wnList_res_re_rawIn_43_sExp[2:0],10'h331}; // @[Cat.scala 33:92]
  wire [16:0] _wnList_res_re_T_375 = {1'h0,wnList_res_re_rawIn_43_sExp[5:3],wnList_res_re_rawIn_43_sExp[2:0],10'h2d7}; // @[Cat.scala 33:92]
  wire [16:0] _wnList_res_re_T_383 = {1'h0,wnList_res_re_rawIn_43_sExp[5:3],wnList_res_re_rawIn_43_sExp[2:0],10'h27b}; // @[Cat.scala 33:92]
  wire [16:0] _wnList_res_re_T_391 = {1'h0,wnList_res_re_rawIn_43_sExp[5:3],wnList_res_re_rawIn_43_sExp[2:0],10'h21f}; // @[Cat.scala 33:92]
  wire [16:0] _wnList_res_re_T_399 = {1'h0,wnList_res_re_rawIn_43_sExp[5:3],wnList_res_re_rawIn_43_sExp[2:0],10'h1c2}; // @[Cat.scala 33:92]
  wire [16:0] _wnList_res_re_T_407 = {1'h0,wnList_res_re_rawIn_43_sExp[5:3],wnList_res_re_rawIn_43_sExp[2:0],10'h163}; // @[Cat.scala 33:92]
  wire [16:0] _wnList_res_re_T_415 = {1'h0,wnList_res_re_rawIn_43_sExp[5:3],wnList_res_re_rawIn_43_sExp[2:0],10'h104}; // @[Cat.scala 33:92]
  wire [16:0] _wnList_res_re_T_423 = {1'h0,wnList_res_re_rawIn_43_sExp[5:3],wnList_res_re_rawIn_43_sExp[2:0],10'ha5}; // @[Cat.scala 33:92]
  wire [16:0] _wnList_res_re_T_431 = {1'h0,wnList_res_re_rawIn_43_sExp[5:3],wnList_res_re_rawIn_43_sExp[2:0],10'h44}; // @[Cat.scala 33:92]
  wire [6:0] wnList_res_re_rawIn_54_sExp = {1'b0,$signed(6'h1d)}; // @[rawFloatFromFN.scala 70:48]
  wire [16:0] _wnList_res_re_T_439 = {1'h0,wnList_res_re_rawIn_54_sExp[5:3],wnList_res_re_rawIn_54_sExp[2:0],10'h3c6}; // @[Cat.scala 33:92]
  wire [16:0] _wnList_res_re_T_447 = {1'h0,wnList_res_re_rawIn_54_sExp[5:3],wnList_res_re_rawIn_54_sExp[2:0],10'h302}; // @[Cat.scala 33:92]
  wire [16:0] _wnList_res_re_T_455 = {1'h0,wnList_res_re_rawIn_54_sExp[5:3],wnList_res_re_rawIn_54_sExp[2:0],10'h23e}; // @[Cat.scala 33:92]
  wire [16:0] _wnList_res_re_T_463 = {1'h0,wnList_res_re_rawIn_54_sExp[5:3],wnList_res_re_rawIn_54_sExp[2:0],10'h178}; // @[Cat.scala 33:92]
  wire [16:0] _wnList_res_re_T_471 = {1'h0,wnList_res_re_rawIn_54_sExp[5:3],wnList_res_re_rawIn_54_sExp[2:0],10'hb2}; // @[Cat.scala 33:92]
  wire [6:0] wnList_res_re_rawIn_59_sExp = {1'b0,$signed(6'h1c)}; // @[rawFloatFromFN.scala 70:48]
  wire [16:0] _wnList_res_re_T_479 = {1'h0,wnList_res_re_rawIn_59_sExp[5:3],wnList_res_re_rawIn_59_sExp[2:0],10'h3d5}; // @[Cat.scala 33:92]
  wire [16:0] _wnList_res_re_T_487 = {1'h0,wnList_res_re_rawIn_59_sExp[5:3],wnList_res_re_rawIn_59_sExp[2:0],10'h245}; // @[Cat.scala 33:92]
  wire [16:0] _wnList_res_re_T_495 = {1'h0,wnList_res_re_rawIn_59_sExp[5:3],wnList_res_re_rawIn_59_sExp[2:0],10'hb5}; // @[Cat.scala 33:92]
  wire [6:0] wnList_res_re_rawIn_62_sExp = {1'b0,$signed(6'h1b)}; // @[rawFloatFromFN.scala 70:48]
  wire [16:0] _wnList_res_re_T_503 = {1'h0,wnList_res_re_rawIn_62_sExp[5:3],wnList_res_re_rawIn_62_sExp[2:0],10'h247}; // @[Cat.scala 33:92]
  wire [6:0] wnList_res_re_rawIn_63_sExp = {1'b0,$signed(6'h1a)}; // @[rawFloatFromFN.scala 70:48]
  wire [16:0] _wnList_res_re_T_511 = {1'h0,wnList_res_re_rawIn_63_sExp[5:3],wnList_res_re_rawIn_63_sExp[2:0],10'h248}; // @[Cat.scala 33:92]
  wire [6:0] wnList_res_re_rawIn_64_sExp = {1'b0,$signed(6'h8)}; // @[rawFloatFromFN.scala 70:48]
  wire [16:0] _wnList_res_re_T_519 = {4'h0,wnList_res_re_rawIn_64_sExp[2:0],10'h0}; // @[Cat.scala 33:92]
  wire [16:0] _wnList_res_re_T_527 = {1'h1,wnList_res_re_rawIn_63_sExp[5:3],wnList_res_re_rawIn_63_sExp[2:0],10'h248}; // @[Cat.scala 33:92]
  wire [16:0] _wnList_res_re_T_535 = {1'h1,wnList_res_re_rawIn_62_sExp[5:3],wnList_res_re_rawIn_62_sExp[2:0],10'h247}; // @[Cat.scala 33:92]
  wire [16:0] _wnList_res_re_T_543 = {1'h1,wnList_res_re_rawIn_59_sExp[5:3],wnList_res_re_rawIn_59_sExp[2:0],10'hb5}; // @[Cat.scala 33:92]
  wire [16:0] _wnList_res_re_T_551 = {1'h1,wnList_res_re_rawIn_59_sExp[5:3],wnList_res_re_rawIn_59_sExp[2:0],10'h245}; // @[Cat.scala 33:92]
  wire [16:0] _wnList_res_re_T_559 = {1'h1,wnList_res_re_rawIn_59_sExp[5:3],wnList_res_re_rawIn_59_sExp[2:0],10'h3d5}; // @[Cat.scala 33:92]
  wire [16:0] _wnList_res_re_T_567 = {1'h1,wnList_res_re_rawIn_54_sExp[5:3],wnList_res_re_rawIn_54_sExp[2:0],10'hb2}; // @[Cat.scala 33:92]
  wire [16:0] _wnList_res_re_T_575 = {1'h1,wnList_res_re_rawIn_54_sExp[5:3],wnList_res_re_rawIn_54_sExp[2:0],10'h178}; // @[Cat.scala 33:92]
  wire [16:0] _wnList_res_re_T_583 = {1'h1,wnList_res_re_rawIn_54_sExp[5:3],wnList_res_re_rawIn_54_sExp[2:0],10'h23e}; // @[Cat.scala 33:92]
  wire [16:0] _wnList_res_re_T_591 = {1'h1,wnList_res_re_rawIn_54_sExp[5:3],wnList_res_re_rawIn_54_sExp[2:0],10'h302}; // @[Cat.scala 33:92]
  wire [16:0] _wnList_res_re_T_599 = {1'h1,wnList_res_re_rawIn_54_sExp[5:3],wnList_res_re_rawIn_54_sExp[2:0],10'h3c6}; // @[Cat.scala 33:92]
  wire [16:0] _wnList_res_re_T_607 = {1'h1,wnList_res_re_rawIn_43_sExp[5:3],wnList_res_re_rawIn_43_sExp[2:0],10'h44}; // @[Cat.scala 33:92]
  wire [16:0] _wnList_res_re_T_615 = {1'h1,wnList_res_re_rawIn_43_sExp[5:3],wnList_res_re_rawIn_43_sExp[2:0],10'ha5}; // @[Cat.scala 33:92]
  wire [16:0] _wnList_res_re_T_623 = {1'h1,wnList_res_re_rawIn_43_sExp[5:3],wnList_res_re_rawIn_43_sExp[2:0],10'h104}; // @[Cat.scala 33:92]
  wire [16:0] _wnList_res_re_T_631 = {1'h1,wnList_res_re_rawIn_43_sExp[5:3],wnList_res_re_rawIn_43_sExp[2:0],10'h163}; // @[Cat.scala 33:92]
  wire [16:0] _wnList_res_re_T_639 = {1'h1,wnList_res_re_rawIn_43_sExp[5:3],wnList_res_re_rawIn_43_sExp[2:0],10'h1c2}; // @[Cat.scala 33:92]
  wire [16:0] _wnList_res_re_T_647 = {1'h1,wnList_res_re_rawIn_43_sExp[5:3],wnList_res_re_rawIn_43_sExp[2:0],10'h21f}; // @[Cat.scala 33:92]
  wire [16:0] _wnList_res_re_T_655 = {1'h1,wnList_res_re_rawIn_43_sExp[5:3],wnList_res_re_rawIn_43_sExp[2:0],10'h27b}; // @[Cat.scala 33:92]
  wire [16:0] _wnList_res_re_T_663 = {1'h1,wnList_res_re_rawIn_43_sExp[5:3],wnList_res_re_rawIn_43_sExp[2:0],10'h2d7}; // @[Cat.scala 33:92]
  wire [16:0] _wnList_res_re_T_671 = {1'h1,wnList_res_re_rawIn_43_sExp[5:3],wnList_res_re_rawIn_43_sExp[2:0],10'h331}; // @[Cat.scala 33:92]
  wire [16:0] _wnList_res_re_T_679 = {1'h1,wnList_res_re_rawIn_43_sExp[5:3],wnList_res_re_rawIn_43_sExp[2:0],10'h38a}; // @[Cat.scala 33:92]
  wire [16:0] _wnList_res_re_T_687 = {1'h1,wnList_res_re_rawIn_43_sExp[5:3],wnList_res_re_rawIn_43_sExp[2:0],10'h3e2}; // @[Cat.scala 33:92]
  wire [16:0] _wnList_res_re_T_695 = {1'h1,wnList_res_re_rawIn_1_sExp[5:3],wnList_res_re_rawIn_1_sExp[2:0],10'h1c}; // @[Cat.scala 33:92]
  wire [16:0] _wnList_res_re_T_703 = {1'h1,wnList_res_re_rawIn_1_sExp[5:3],wnList_res_re_rawIn_1_sExp[2:0],10'h47}; // @[Cat.scala 33:92]
  wire [16:0] _wnList_res_re_T_711 = {1'h1,wnList_res_re_rawIn_1_sExp[5:3],wnList_res_re_rawIn_1_sExp[2:0],10'h71}; // @[Cat.scala 33:92]
  wire [16:0] _wnList_res_re_T_719 = {1'h1,wnList_res_re_rawIn_1_sExp[5:3],wnList_res_re_rawIn_1_sExp[2:0],10'h9b}; // @[Cat.scala 33:92]
  wire [16:0] _wnList_res_re_T_727 = {1'h1,wnList_res_re_rawIn_1_sExp[5:3],wnList_res_re_rawIn_1_sExp[2:0],10'hc3}; // @[Cat.scala 33:92]
  wire [16:0] _wnList_res_re_T_735 = {1'h1,wnList_res_re_rawIn_1_sExp[5:3],wnList_res_re_rawIn_1_sExp[2:0],10'heb}; // @[Cat.scala 33:92]
  wire [16:0] _wnList_res_re_T_743 = {1'h1,wnList_res_re_rawIn_1_sExp[5:3],wnList_res_re_rawIn_1_sExp[2:0],10'h113}; // @[Cat.scala 33:92]
  wire [16:0] _wnList_res_re_T_751 = {1'h1,wnList_res_re_rawIn_1_sExp[5:3],wnList_res_re_rawIn_1_sExp[2:0],10'h139}; // @[Cat.scala 33:92]
  wire [16:0] _wnList_res_re_T_759 = {1'h1,wnList_res_re_rawIn_1_sExp[5:3],wnList_res_re_rawIn_1_sExp[2:0],10'h15f}; // @[Cat.scala 33:92]
  wire [16:0] _wnList_res_re_T_767 = {1'h1,wnList_res_re_rawIn_1_sExp[5:3],wnList_res_re_rawIn_1_sExp[2:0],10'h184}; // @[Cat.scala 33:92]
  wire [16:0] _wnList_res_re_T_775 = {1'h1,wnList_res_re_rawIn_1_sExp[5:3],wnList_res_re_rawIn_1_sExp[2:0],10'h1a8}; // @[Cat.scala 33:92]
  wire [16:0] _wnList_res_re_T_783 = {1'h1,wnList_res_re_rawIn_1_sExp[5:3],wnList_res_re_rawIn_1_sExp[2:0],10'h1cb}; // @[Cat.scala 33:92]
  wire [16:0] _wnList_res_re_T_791 = {1'h1,wnList_res_re_rawIn_1_sExp[5:3],wnList_res_re_rawIn_1_sExp[2:0],10'h1ed}; // @[Cat.scala 33:92]
  wire [16:0] _wnList_res_re_T_799 = {1'h1,wnList_res_re_rawIn_1_sExp[5:3],wnList_res_re_rawIn_1_sExp[2:0],10'h20e}; // @[Cat.scala 33:92]
  wire [16:0] _wnList_res_re_T_807 = {1'h1,wnList_res_re_rawIn_1_sExp[5:3],wnList_res_re_rawIn_1_sExp[2:0],10'h22f}; // @[Cat.scala 33:92]
  wire [16:0] _wnList_res_re_T_815 = {1'h1,wnList_res_re_rawIn_1_sExp[5:3],wnList_res_re_rawIn_1_sExp[2:0],10'h24e}; // @[Cat.scala 33:92]
  wire [16:0] _wnList_res_re_T_823 = {1'h1,wnList_res_re_rawIn_1_sExp[5:3],wnList_res_re_rawIn_1_sExp[2:0],10'h26c}; // @[Cat.scala 33:92]
  wire [16:0] _wnList_res_re_T_831 = {1'h1,wnList_res_re_rawIn_1_sExp[5:3],wnList_res_re_rawIn_1_sExp[2:0],10'h28a}; // @[Cat.scala 33:92]
  wire [16:0] _wnList_res_re_T_839 = {1'h1,wnList_res_re_rawIn_1_sExp[5:3],wnList_res_re_rawIn_1_sExp[2:0],10'h2a6}; // @[Cat.scala 33:92]
  wire [16:0] _wnList_res_re_T_847 = {1'h1,wnList_res_re_rawIn_1_sExp[5:3],wnList_res_re_rawIn_1_sExp[2:0],10'h2c2}; // @[Cat.scala 33:92]
  wire [16:0] _wnList_res_re_T_855 = {1'h1,wnList_res_re_rawIn_1_sExp[5:3],wnList_res_re_rawIn_1_sExp[2:0],10'h2dc}; // @[Cat.scala 33:92]
  wire [16:0] _wnList_res_re_T_863 = {1'h1,wnList_res_re_rawIn_1_sExp[5:3],wnList_res_re_rawIn_1_sExp[2:0],10'h2f5}; // @[Cat.scala 33:92]
  wire [16:0] _wnList_res_re_T_871 = {1'h1,wnList_res_re_rawIn_1_sExp[5:3],wnList_res_re_rawIn_1_sExp[2:0],10'h30e}; // @[Cat.scala 33:92]
  wire [16:0] _wnList_res_re_T_879 = {1'h1,wnList_res_re_rawIn_1_sExp[5:3],wnList_res_re_rawIn_1_sExp[2:0],10'h325}; // @[Cat.scala 33:92]
  wire [16:0] _wnList_res_re_T_887 = {1'h1,wnList_res_re_rawIn_1_sExp[5:3],wnList_res_re_rawIn_1_sExp[2:0],10'h33b}; // @[Cat.scala 33:92]
  wire [16:0] _wnList_res_re_T_895 = {1'h1,wnList_res_re_rawIn_1_sExp[5:3],wnList_res_re_rawIn_1_sExp[2:0],10'h350}; // @[Cat.scala 33:92]
  wire [16:0] _wnList_res_re_T_903 = {1'h1,wnList_res_re_rawIn_1_sExp[5:3],wnList_res_re_rawIn_1_sExp[2:0],10'h364}; // @[Cat.scala 33:92]
  wire [16:0] _wnList_res_re_T_911 = {1'h1,wnList_res_re_rawIn_1_sExp[5:3],wnList_res_re_rawIn_1_sExp[2:0],10'h376}; // @[Cat.scala 33:92]
  wire [16:0] _wnList_res_re_T_919 = {1'h1,wnList_res_re_rawIn_1_sExp[5:3],wnList_res_re_rawIn_1_sExp[2:0],10'h388}; // @[Cat.scala 33:92]
  wire [16:0] _wnList_res_re_T_927 = {1'h1,wnList_res_re_rawIn_1_sExp[5:3],wnList_res_re_rawIn_1_sExp[2:0],10'h398}; // @[Cat.scala 33:92]
  wire [16:0] _wnList_res_re_T_935 = {1'h1,wnList_res_re_rawIn_1_sExp[5:3],wnList_res_re_rawIn_1_sExp[2:0],10'h3a7}; // @[Cat.scala 33:92]
  wire [16:0] _wnList_res_re_T_943 = {1'h1,wnList_res_re_rawIn_1_sExp[5:3],wnList_res_re_rawIn_1_sExp[2:0],10'h3b5}; // @[Cat.scala 33:92]
  wire [16:0] _wnList_res_re_T_951 = {1'h1,wnList_res_re_rawIn_1_sExp[5:3],wnList_res_re_rawIn_1_sExp[2:0],10'h3c2}; // @[Cat.scala 33:92]
  wire [16:0] _wnList_res_re_T_959 = {1'h1,wnList_res_re_rawIn_1_sExp[5:3],wnList_res_re_rawIn_1_sExp[2:0],10'h3ce}; // @[Cat.scala 33:92]
  wire [16:0] _wnList_res_re_T_967 = {1'h1,wnList_res_re_rawIn_1_sExp[5:3],wnList_res_re_rawIn_1_sExp[2:0],10'h3d8}; // @[Cat.scala 33:92]
  wire [16:0] _wnList_res_re_T_975 = {1'h1,wnList_res_re_rawIn_1_sExp[5:3],wnList_res_re_rawIn_1_sExp[2:0],10'h3e1}; // @[Cat.scala 33:92]
  wire [16:0] _wnList_res_re_T_983 = {1'h1,wnList_res_re_rawIn_1_sExp[5:3],wnList_res_re_rawIn_1_sExp[2:0],10'h3e9}; // @[Cat.scala 33:92]
  wire [16:0] _wnList_res_re_T_991 = {1'h1,wnList_res_re_rawIn_1_sExp[5:3],wnList_res_re_rawIn_1_sExp[2:0],10'h3f0}; // @[Cat.scala 33:92]
  wire [16:0] _wnList_res_re_T_999 = {1'h1,wnList_res_re_rawIn_1_sExp[5:3],wnList_res_re_rawIn_1_sExp[2:0],10'h3f6}; // @[Cat.scala 33:92]
  wire [16:0] _wnList_res_re_T_1007 = {1'h1,wnList_res_re_rawIn_1_sExp[5:3],wnList_res_re_rawIn_1_sExp[2:0],10'h3fa}; // @[Cat.scala 33:92]
  wire [16:0] _wnList_res_re_T_1015 = {1'h1,wnList_res_re_rawIn_1_sExp[5:3],wnList_res_re_rawIn_1_sExp[2:0],10'h3fd}; // @[Cat.scala 33:92]
  wire [16:0] _wnList_res_re_T_1023 = {1'h1,wnList_res_re_rawIn_1_sExp[5:3],wnList_res_re_rawIn_1_sExp[2:0],10'h3ff}; // @[Cat.scala 33:92]
  wire [16:0] _GEN_2 = 7'h1 == _wnList_T[6:0] ? _wnList_res_re_T_15 : _wnList_res_re_T_7; // @[FFT.scala 104:{12,12}]
  wire [16:0] _GEN_3 = 7'h2 == _wnList_T[6:0] ? _wnList_res_re_T_23 : _GEN_2; // @[FFT.scala 104:{12,12}]
  wire [16:0] _GEN_4 = 7'h3 == _wnList_T[6:0] ? _wnList_res_re_T_31 : _GEN_3; // @[FFT.scala 104:{12,12}]
  wire [16:0] _GEN_5 = 7'h4 == _wnList_T[6:0] ? _wnList_res_re_T_39 : _GEN_4; // @[FFT.scala 104:{12,12}]
  wire [16:0] _GEN_6 = 7'h5 == _wnList_T[6:0] ? _wnList_res_re_T_47 : _GEN_5; // @[FFT.scala 104:{12,12}]
  wire [16:0] _GEN_7 = 7'h6 == _wnList_T[6:0] ? _wnList_res_re_T_55 : _GEN_6; // @[FFT.scala 104:{12,12}]
  wire [16:0] _GEN_8 = 7'h7 == _wnList_T[6:0] ? _wnList_res_re_T_63 : _GEN_7; // @[FFT.scala 104:{12,12}]
  wire [16:0] _GEN_9 = 7'h8 == _wnList_T[6:0] ? _wnList_res_re_T_71 : _GEN_8; // @[FFT.scala 104:{12,12}]
  wire [16:0] _GEN_10 = 7'h9 == _wnList_T[6:0] ? _wnList_res_re_T_79 : _GEN_9; // @[FFT.scala 104:{12,12}]
  wire [16:0] _GEN_11 = 7'ha == _wnList_T[6:0] ? _wnList_res_re_T_87 : _GEN_10; // @[FFT.scala 104:{12,12}]
  wire [16:0] _GEN_12 = 7'hb == _wnList_T[6:0] ? _wnList_res_re_T_95 : _GEN_11; // @[FFT.scala 104:{12,12}]
  wire [16:0] _GEN_13 = 7'hc == _wnList_T[6:0] ? _wnList_res_re_T_103 : _GEN_12; // @[FFT.scala 104:{12,12}]
  wire [16:0] _GEN_14 = 7'hd == _wnList_T[6:0] ? _wnList_res_re_T_111 : _GEN_13; // @[FFT.scala 104:{12,12}]
  wire [16:0] _GEN_15 = 7'he == _wnList_T[6:0] ? _wnList_res_re_T_119 : _GEN_14; // @[FFT.scala 104:{12,12}]
  wire [16:0] _GEN_16 = 7'hf == _wnList_T[6:0] ? _wnList_res_re_T_127 : _GEN_15; // @[FFT.scala 104:{12,12}]
  wire [16:0] _GEN_17 = 7'h10 == _wnList_T[6:0] ? _wnList_res_re_T_135 : _GEN_16; // @[FFT.scala 104:{12,12}]
  wire [16:0] _GEN_18 = 7'h11 == _wnList_T[6:0] ? _wnList_res_re_T_143 : _GEN_17; // @[FFT.scala 104:{12,12}]
  wire [16:0] _GEN_19 = 7'h12 == _wnList_T[6:0] ? _wnList_res_re_T_151 : _GEN_18; // @[FFT.scala 104:{12,12}]
  wire [16:0] _GEN_20 = 7'h13 == _wnList_T[6:0] ? _wnList_res_re_T_159 : _GEN_19; // @[FFT.scala 104:{12,12}]
  wire [16:0] _GEN_21 = 7'h14 == _wnList_T[6:0] ? _wnList_res_re_T_167 : _GEN_20; // @[FFT.scala 104:{12,12}]
  wire [16:0] _GEN_22 = 7'h15 == _wnList_T[6:0] ? _wnList_res_re_T_175 : _GEN_21; // @[FFT.scala 104:{12,12}]
  wire [16:0] _GEN_23 = 7'h16 == _wnList_T[6:0] ? _wnList_res_re_T_183 : _GEN_22; // @[FFT.scala 104:{12,12}]
  wire [16:0] _GEN_24 = 7'h17 == _wnList_T[6:0] ? _wnList_res_re_T_191 : _GEN_23; // @[FFT.scala 104:{12,12}]
  wire [16:0] _GEN_25 = 7'h18 == _wnList_T[6:0] ? _wnList_res_re_T_199 : _GEN_24; // @[FFT.scala 104:{12,12}]
  wire [16:0] _GEN_26 = 7'h19 == _wnList_T[6:0] ? _wnList_res_re_T_207 : _GEN_25; // @[FFT.scala 104:{12,12}]
  wire [16:0] _GEN_27 = 7'h1a == _wnList_T[6:0] ? _wnList_res_re_T_215 : _GEN_26; // @[FFT.scala 104:{12,12}]
  wire [16:0] _GEN_28 = 7'h1b == _wnList_T[6:0] ? _wnList_res_re_T_223 : _GEN_27; // @[FFT.scala 104:{12,12}]
  wire [16:0] _GEN_29 = 7'h1c == _wnList_T[6:0] ? _wnList_res_re_T_231 : _GEN_28; // @[FFT.scala 104:{12,12}]
  wire [16:0] _GEN_30 = 7'h1d == _wnList_T[6:0] ? _wnList_res_re_T_239 : _GEN_29; // @[FFT.scala 104:{12,12}]
  wire [16:0] _GEN_31 = 7'h1e == _wnList_T[6:0] ? _wnList_res_re_T_247 : _GEN_30; // @[FFT.scala 104:{12,12}]
  wire [16:0] _GEN_32 = 7'h1f == _wnList_T[6:0] ? _wnList_res_re_T_255 : _GEN_31; // @[FFT.scala 104:{12,12}]
  wire [16:0] _GEN_33 = 7'h20 == _wnList_T[6:0] ? _wnList_res_re_T_263 : _GEN_32; // @[FFT.scala 104:{12,12}]
  wire [16:0] _GEN_34 = 7'h21 == _wnList_T[6:0] ? _wnList_res_re_T_271 : _GEN_33; // @[FFT.scala 104:{12,12}]
  wire [16:0] _GEN_35 = 7'h22 == _wnList_T[6:0] ? _wnList_res_re_T_279 : _GEN_34; // @[FFT.scala 104:{12,12}]
  wire [16:0] _GEN_36 = 7'h23 == _wnList_T[6:0] ? _wnList_res_re_T_287 : _GEN_35; // @[FFT.scala 104:{12,12}]
  wire [16:0] _GEN_37 = 7'h24 == _wnList_T[6:0] ? _wnList_res_re_T_295 : _GEN_36; // @[FFT.scala 104:{12,12}]
  wire [16:0] _GEN_38 = 7'h25 == _wnList_T[6:0] ? _wnList_res_re_T_303 : _GEN_37; // @[FFT.scala 104:{12,12}]
  wire [16:0] _GEN_39 = 7'h26 == _wnList_T[6:0] ? _wnList_res_re_T_311 : _GEN_38; // @[FFT.scala 104:{12,12}]
  wire [16:0] _GEN_40 = 7'h27 == _wnList_T[6:0] ? _wnList_res_re_T_319 : _GEN_39; // @[FFT.scala 104:{12,12}]
  wire [16:0] _GEN_41 = 7'h28 == _wnList_T[6:0] ? _wnList_res_re_T_327 : _GEN_40; // @[FFT.scala 104:{12,12}]
  wire [16:0] _GEN_42 = 7'h29 == _wnList_T[6:0] ? _wnList_res_re_T_335 : _GEN_41; // @[FFT.scala 104:{12,12}]
  wire [16:0] _GEN_43 = 7'h2a == _wnList_T[6:0] ? _wnList_res_re_T_343 : _GEN_42; // @[FFT.scala 104:{12,12}]
  wire [16:0] _GEN_44 = 7'h2b == _wnList_T[6:0] ? _wnList_res_re_T_351 : _GEN_43; // @[FFT.scala 104:{12,12}]
  wire [16:0] _GEN_45 = 7'h2c == _wnList_T[6:0] ? _wnList_res_re_T_359 : _GEN_44; // @[FFT.scala 104:{12,12}]
  wire [16:0] _GEN_46 = 7'h2d == _wnList_T[6:0] ? _wnList_res_re_T_367 : _GEN_45; // @[FFT.scala 104:{12,12}]
  wire [16:0] _GEN_47 = 7'h2e == _wnList_T[6:0] ? _wnList_res_re_T_375 : _GEN_46; // @[FFT.scala 104:{12,12}]
  wire [16:0] _GEN_48 = 7'h2f == _wnList_T[6:0] ? _wnList_res_re_T_383 : _GEN_47; // @[FFT.scala 104:{12,12}]
  wire [16:0] _GEN_49 = 7'h30 == _wnList_T[6:0] ? _wnList_res_re_T_391 : _GEN_48; // @[FFT.scala 104:{12,12}]
  wire [16:0] _GEN_50 = 7'h31 == _wnList_T[6:0] ? _wnList_res_re_T_399 : _GEN_49; // @[FFT.scala 104:{12,12}]
  wire [16:0] _GEN_51 = 7'h32 == _wnList_T[6:0] ? _wnList_res_re_T_407 : _GEN_50; // @[FFT.scala 104:{12,12}]
  wire [16:0] _GEN_52 = 7'h33 == _wnList_T[6:0] ? _wnList_res_re_T_415 : _GEN_51; // @[FFT.scala 104:{12,12}]
  wire [16:0] _GEN_53 = 7'h34 == _wnList_T[6:0] ? _wnList_res_re_T_423 : _GEN_52; // @[FFT.scala 104:{12,12}]
  wire [16:0] _GEN_54 = 7'h35 == _wnList_T[6:0] ? _wnList_res_re_T_431 : _GEN_53; // @[FFT.scala 104:{12,12}]
  wire [16:0] _GEN_55 = 7'h36 == _wnList_T[6:0] ? _wnList_res_re_T_439 : _GEN_54; // @[FFT.scala 104:{12,12}]
  wire [16:0] _GEN_56 = 7'h37 == _wnList_T[6:0] ? _wnList_res_re_T_447 : _GEN_55; // @[FFT.scala 104:{12,12}]
  wire [16:0] _GEN_57 = 7'h38 == _wnList_T[6:0] ? _wnList_res_re_T_455 : _GEN_56; // @[FFT.scala 104:{12,12}]
  wire [16:0] _GEN_58 = 7'h39 == _wnList_T[6:0] ? _wnList_res_re_T_463 : _GEN_57; // @[FFT.scala 104:{12,12}]
  wire [16:0] _GEN_59 = 7'h3a == _wnList_T[6:0] ? _wnList_res_re_T_471 : _GEN_58; // @[FFT.scala 104:{12,12}]
  wire [16:0] _GEN_60 = 7'h3b == _wnList_T[6:0] ? _wnList_res_re_T_479 : _GEN_59; // @[FFT.scala 104:{12,12}]
  wire [16:0] _GEN_61 = 7'h3c == _wnList_T[6:0] ? _wnList_res_re_T_487 : _GEN_60; // @[FFT.scala 104:{12,12}]
  wire [16:0] _GEN_62 = 7'h3d == _wnList_T[6:0] ? _wnList_res_re_T_495 : _GEN_61; // @[FFT.scala 104:{12,12}]
  wire [16:0] _GEN_63 = 7'h3e == _wnList_T[6:0] ? _wnList_res_re_T_503 : _GEN_62; // @[FFT.scala 104:{12,12}]
  wire [16:0] _GEN_64 = 7'h3f == _wnList_T[6:0] ? _wnList_res_re_T_511 : _GEN_63; // @[FFT.scala 104:{12,12}]
  wire [16:0] _GEN_65 = 7'h40 == _wnList_T[6:0] ? _wnList_res_re_T_519 : _GEN_64; // @[FFT.scala 104:{12,12}]
  wire [16:0] _GEN_66 = 7'h41 == _wnList_T[6:0] ? _wnList_res_re_T_527 : _GEN_65; // @[FFT.scala 104:{12,12}]
  wire [16:0] _GEN_67 = 7'h42 == _wnList_T[6:0] ? _wnList_res_re_T_535 : _GEN_66; // @[FFT.scala 104:{12,12}]
  wire [16:0] _GEN_68 = 7'h43 == _wnList_T[6:0] ? _wnList_res_re_T_543 : _GEN_67; // @[FFT.scala 104:{12,12}]
  wire [16:0] _GEN_69 = 7'h44 == _wnList_T[6:0] ? _wnList_res_re_T_551 : _GEN_68; // @[FFT.scala 104:{12,12}]
  wire [16:0] _GEN_70 = 7'h45 == _wnList_T[6:0] ? _wnList_res_re_T_559 : _GEN_69; // @[FFT.scala 104:{12,12}]
  wire [16:0] _GEN_71 = 7'h46 == _wnList_T[6:0] ? _wnList_res_re_T_567 : _GEN_70; // @[FFT.scala 104:{12,12}]
  wire [16:0] _GEN_72 = 7'h47 == _wnList_T[6:0] ? _wnList_res_re_T_575 : _GEN_71; // @[FFT.scala 104:{12,12}]
  wire [16:0] _GEN_73 = 7'h48 == _wnList_T[6:0] ? _wnList_res_re_T_583 : _GEN_72; // @[FFT.scala 104:{12,12}]
  wire [16:0] _GEN_74 = 7'h49 == _wnList_T[6:0] ? _wnList_res_re_T_591 : _GEN_73; // @[FFT.scala 104:{12,12}]
  wire [16:0] _GEN_75 = 7'h4a == _wnList_T[6:0] ? _wnList_res_re_T_599 : _GEN_74; // @[FFT.scala 104:{12,12}]
  wire [16:0] _GEN_76 = 7'h4b == _wnList_T[6:0] ? _wnList_res_re_T_607 : _GEN_75; // @[FFT.scala 104:{12,12}]
  wire [16:0] _GEN_77 = 7'h4c == _wnList_T[6:0] ? _wnList_res_re_T_615 : _GEN_76; // @[FFT.scala 104:{12,12}]
  wire [16:0] _GEN_78 = 7'h4d == _wnList_T[6:0] ? _wnList_res_re_T_623 : _GEN_77; // @[FFT.scala 104:{12,12}]
  wire [16:0] _GEN_79 = 7'h4e == _wnList_T[6:0] ? _wnList_res_re_T_631 : _GEN_78; // @[FFT.scala 104:{12,12}]
  wire [16:0] _GEN_80 = 7'h4f == _wnList_T[6:0] ? _wnList_res_re_T_639 : _GEN_79; // @[FFT.scala 104:{12,12}]
  wire [16:0] _GEN_81 = 7'h50 == _wnList_T[6:0] ? _wnList_res_re_T_647 : _GEN_80; // @[FFT.scala 104:{12,12}]
  wire [16:0] _GEN_82 = 7'h51 == _wnList_T[6:0] ? _wnList_res_re_T_655 : _GEN_81; // @[FFT.scala 104:{12,12}]
  wire [16:0] _GEN_83 = 7'h52 == _wnList_T[6:0] ? _wnList_res_re_T_663 : _GEN_82; // @[FFT.scala 104:{12,12}]
  wire [16:0] _GEN_84 = 7'h53 == _wnList_T[6:0] ? _wnList_res_re_T_671 : _GEN_83; // @[FFT.scala 104:{12,12}]
  wire [16:0] _GEN_85 = 7'h54 == _wnList_T[6:0] ? _wnList_res_re_T_679 : _GEN_84; // @[FFT.scala 104:{12,12}]
  wire [16:0] _GEN_86 = 7'h55 == _wnList_T[6:0] ? _wnList_res_re_T_687 : _GEN_85; // @[FFT.scala 104:{12,12}]
  wire [16:0] _GEN_87 = 7'h56 == _wnList_T[6:0] ? _wnList_res_re_T_695 : _GEN_86; // @[FFT.scala 104:{12,12}]
  wire [16:0] _GEN_88 = 7'h57 == _wnList_T[6:0] ? _wnList_res_re_T_703 : _GEN_87; // @[FFT.scala 104:{12,12}]
  wire [16:0] _GEN_89 = 7'h58 == _wnList_T[6:0] ? _wnList_res_re_T_711 : _GEN_88; // @[FFT.scala 104:{12,12}]
  wire [16:0] _GEN_90 = 7'h59 == _wnList_T[6:0] ? _wnList_res_re_T_719 : _GEN_89; // @[FFT.scala 104:{12,12}]
  wire [16:0] _GEN_91 = 7'h5a == _wnList_T[6:0] ? _wnList_res_re_T_727 : _GEN_90; // @[FFT.scala 104:{12,12}]
  wire [16:0] _GEN_92 = 7'h5b == _wnList_T[6:0] ? _wnList_res_re_T_735 : _GEN_91; // @[FFT.scala 104:{12,12}]
  wire [16:0] _GEN_93 = 7'h5c == _wnList_T[6:0] ? _wnList_res_re_T_743 : _GEN_92; // @[FFT.scala 104:{12,12}]
  wire [16:0] _GEN_94 = 7'h5d == _wnList_T[6:0] ? _wnList_res_re_T_751 : _GEN_93; // @[FFT.scala 104:{12,12}]
  wire [16:0] _GEN_95 = 7'h5e == _wnList_T[6:0] ? _wnList_res_re_T_759 : _GEN_94; // @[FFT.scala 104:{12,12}]
  wire [16:0] _GEN_96 = 7'h5f == _wnList_T[6:0] ? _wnList_res_re_T_767 : _GEN_95; // @[FFT.scala 104:{12,12}]
  wire [16:0] _GEN_97 = 7'h60 == _wnList_T[6:0] ? _wnList_res_re_T_775 : _GEN_96; // @[FFT.scala 104:{12,12}]
  wire [16:0] _GEN_98 = 7'h61 == _wnList_T[6:0] ? _wnList_res_re_T_783 : _GEN_97; // @[FFT.scala 104:{12,12}]
  wire [16:0] _GEN_99 = 7'h62 == _wnList_T[6:0] ? _wnList_res_re_T_791 : _GEN_98; // @[FFT.scala 104:{12,12}]
  wire [16:0] _GEN_100 = 7'h63 == _wnList_T[6:0] ? _wnList_res_re_T_799 : _GEN_99; // @[FFT.scala 104:{12,12}]
  wire [16:0] _GEN_101 = 7'h64 == _wnList_T[6:0] ? _wnList_res_re_T_807 : _GEN_100; // @[FFT.scala 104:{12,12}]
  wire [16:0] _GEN_102 = 7'h65 == _wnList_T[6:0] ? _wnList_res_re_T_815 : _GEN_101; // @[FFT.scala 104:{12,12}]
  wire [16:0] _GEN_103 = 7'h66 == _wnList_T[6:0] ? _wnList_res_re_T_823 : _GEN_102; // @[FFT.scala 104:{12,12}]
  wire [16:0] _GEN_104 = 7'h67 == _wnList_T[6:0] ? _wnList_res_re_T_831 : _GEN_103; // @[FFT.scala 104:{12,12}]
  wire [16:0] _GEN_105 = 7'h68 == _wnList_T[6:0] ? _wnList_res_re_T_839 : _GEN_104; // @[FFT.scala 104:{12,12}]
  wire [16:0] _GEN_106 = 7'h69 == _wnList_T[6:0] ? _wnList_res_re_T_847 : _GEN_105; // @[FFT.scala 104:{12,12}]
  wire [16:0] _GEN_107 = 7'h6a == _wnList_T[6:0] ? _wnList_res_re_T_855 : _GEN_106; // @[FFT.scala 104:{12,12}]
  wire [16:0] _GEN_108 = 7'h6b == _wnList_T[6:0] ? _wnList_res_re_T_863 : _GEN_107; // @[FFT.scala 104:{12,12}]
  wire [16:0] _GEN_109 = 7'h6c == _wnList_T[6:0] ? _wnList_res_re_T_871 : _GEN_108; // @[FFT.scala 104:{12,12}]
  wire [16:0] _GEN_110 = 7'h6d == _wnList_T[6:0] ? _wnList_res_re_T_879 : _GEN_109; // @[FFT.scala 104:{12,12}]
  wire [16:0] _GEN_111 = 7'h6e == _wnList_T[6:0] ? _wnList_res_re_T_887 : _GEN_110; // @[FFT.scala 104:{12,12}]
  wire [16:0] _GEN_112 = 7'h6f == _wnList_T[6:0] ? _wnList_res_re_T_895 : _GEN_111; // @[FFT.scala 104:{12,12}]
  wire [16:0] _GEN_113 = 7'h70 == _wnList_T[6:0] ? _wnList_res_re_T_903 : _GEN_112; // @[FFT.scala 104:{12,12}]
  wire [16:0] _GEN_114 = 7'h71 == _wnList_T[6:0] ? _wnList_res_re_T_911 : _GEN_113; // @[FFT.scala 104:{12,12}]
  wire [16:0] _GEN_115 = 7'h72 == _wnList_T[6:0] ? _wnList_res_re_T_919 : _GEN_114; // @[FFT.scala 104:{12,12}]
  wire [16:0] _GEN_116 = 7'h73 == _wnList_T[6:0] ? _wnList_res_re_T_927 : _GEN_115; // @[FFT.scala 104:{12,12}]
  wire [16:0] _GEN_117 = 7'h74 == _wnList_T[6:0] ? _wnList_res_re_T_935 : _GEN_116; // @[FFT.scala 104:{12,12}]
  wire [16:0] _GEN_118 = 7'h75 == _wnList_T[6:0] ? _wnList_res_re_T_943 : _GEN_117; // @[FFT.scala 104:{12,12}]
  wire [16:0] _GEN_119 = 7'h76 == _wnList_T[6:0] ? _wnList_res_re_T_951 : _GEN_118; // @[FFT.scala 104:{12,12}]
  wire [16:0] _GEN_120 = 7'h77 == _wnList_T[6:0] ? _wnList_res_re_T_959 : _GEN_119; // @[FFT.scala 104:{12,12}]
  wire [16:0] _GEN_121 = 7'h78 == _wnList_T[6:0] ? _wnList_res_re_T_967 : _GEN_120; // @[FFT.scala 104:{12,12}]
  wire [16:0] _GEN_122 = 7'h79 == _wnList_T[6:0] ? _wnList_res_re_T_975 : _GEN_121; // @[FFT.scala 104:{12,12}]
  wire [16:0] _GEN_123 = 7'h7a == _wnList_T[6:0] ? _wnList_res_re_T_983 : _GEN_122; // @[FFT.scala 104:{12,12}]
  wire [16:0] _GEN_124 = 7'h7b == _wnList_T[6:0] ? _wnList_res_re_T_991 : _GEN_123; // @[FFT.scala 104:{12,12}]
  wire [16:0] _GEN_125 = 7'h7c == _wnList_T[6:0] ? _wnList_res_re_T_999 : _GEN_124; // @[FFT.scala 104:{12,12}]
  wire [16:0] _GEN_126 = 7'h7d == _wnList_T[6:0] ? _wnList_res_re_T_1007 : _GEN_125; // @[FFT.scala 104:{12,12}]
  wire [16:0] _GEN_127 = 7'h7e == _wnList_T[6:0] ? _wnList_res_re_T_1015 : _GEN_126; // @[FFT.scala 104:{12,12}]
  wire [16:0] _wnList_res_im_T_519 = {1'h1,wnList_res_re_rawIn__sExp[5:3],wnList_res_re_rawIn__sExp[2:0],10'h0}; // @[Cat.scala 33:92]
  wire [16:0] _GEN_130 = 7'h1 == _wnList_T[6:0] ? _wnList_res_re_T_527 : _wnList_res_re_T_519; // @[FFT.scala 105:{12,12}]
  wire [16:0] _GEN_131 = 7'h2 == _wnList_T[6:0] ? _wnList_res_re_T_535 : _GEN_130; // @[FFT.scala 105:{12,12}]
  wire [16:0] _GEN_132 = 7'h3 == _wnList_T[6:0] ? _wnList_res_re_T_543 : _GEN_131; // @[FFT.scala 105:{12,12}]
  wire [16:0] _GEN_133 = 7'h4 == _wnList_T[6:0] ? _wnList_res_re_T_551 : _GEN_132; // @[FFT.scala 105:{12,12}]
  wire [16:0] _GEN_134 = 7'h5 == _wnList_T[6:0] ? _wnList_res_re_T_559 : _GEN_133; // @[FFT.scala 105:{12,12}]
  wire [16:0] _GEN_135 = 7'h6 == _wnList_T[6:0] ? _wnList_res_re_T_567 : _GEN_134; // @[FFT.scala 105:{12,12}]
  wire [16:0] _GEN_136 = 7'h7 == _wnList_T[6:0] ? _wnList_res_re_T_575 : _GEN_135; // @[FFT.scala 105:{12,12}]
  wire [16:0] _GEN_137 = 7'h8 == _wnList_T[6:0] ? _wnList_res_re_T_583 : _GEN_136; // @[FFT.scala 105:{12,12}]
  wire [16:0] _GEN_138 = 7'h9 == _wnList_T[6:0] ? _wnList_res_re_T_591 : _GEN_137; // @[FFT.scala 105:{12,12}]
  wire [16:0] _GEN_139 = 7'ha == _wnList_T[6:0] ? _wnList_res_re_T_599 : _GEN_138; // @[FFT.scala 105:{12,12}]
  wire [16:0] _GEN_140 = 7'hb == _wnList_T[6:0] ? _wnList_res_re_T_607 : _GEN_139; // @[FFT.scala 105:{12,12}]
  wire [16:0] _GEN_141 = 7'hc == _wnList_T[6:0] ? _wnList_res_re_T_615 : _GEN_140; // @[FFT.scala 105:{12,12}]
  wire [16:0] _GEN_142 = 7'hd == _wnList_T[6:0] ? _wnList_res_re_T_623 : _GEN_141; // @[FFT.scala 105:{12,12}]
  wire [16:0] _GEN_143 = 7'he == _wnList_T[6:0] ? _wnList_res_re_T_631 : _GEN_142; // @[FFT.scala 105:{12,12}]
  wire [16:0] _GEN_144 = 7'hf == _wnList_T[6:0] ? _wnList_res_re_T_639 : _GEN_143; // @[FFT.scala 105:{12,12}]
  wire [16:0] _GEN_145 = 7'h10 == _wnList_T[6:0] ? _wnList_res_re_T_647 : _GEN_144; // @[FFT.scala 105:{12,12}]
  wire [16:0] _GEN_146 = 7'h11 == _wnList_T[6:0] ? _wnList_res_re_T_655 : _GEN_145; // @[FFT.scala 105:{12,12}]
  wire [16:0] _GEN_147 = 7'h12 == _wnList_T[6:0] ? _wnList_res_re_T_663 : _GEN_146; // @[FFT.scala 105:{12,12}]
  wire [16:0] _GEN_148 = 7'h13 == _wnList_T[6:0] ? _wnList_res_re_T_671 : _GEN_147; // @[FFT.scala 105:{12,12}]
  wire [16:0] _GEN_149 = 7'h14 == _wnList_T[6:0] ? _wnList_res_re_T_679 : _GEN_148; // @[FFT.scala 105:{12,12}]
  wire [16:0] _GEN_150 = 7'h15 == _wnList_T[6:0] ? _wnList_res_re_T_687 : _GEN_149; // @[FFT.scala 105:{12,12}]
  wire [16:0] _GEN_151 = 7'h16 == _wnList_T[6:0] ? _wnList_res_re_T_695 : _GEN_150; // @[FFT.scala 105:{12,12}]
  wire [16:0] _GEN_152 = 7'h17 == _wnList_T[6:0] ? _wnList_res_re_T_703 : _GEN_151; // @[FFT.scala 105:{12,12}]
  wire [16:0] _GEN_153 = 7'h18 == _wnList_T[6:0] ? _wnList_res_re_T_711 : _GEN_152; // @[FFT.scala 105:{12,12}]
  wire [16:0] _GEN_154 = 7'h19 == _wnList_T[6:0] ? _wnList_res_re_T_719 : _GEN_153; // @[FFT.scala 105:{12,12}]
  wire [16:0] _GEN_155 = 7'h1a == _wnList_T[6:0] ? _wnList_res_re_T_727 : _GEN_154; // @[FFT.scala 105:{12,12}]
  wire [16:0] _GEN_156 = 7'h1b == _wnList_T[6:0] ? _wnList_res_re_T_735 : _GEN_155; // @[FFT.scala 105:{12,12}]
  wire [16:0] _GEN_157 = 7'h1c == _wnList_T[6:0] ? _wnList_res_re_T_743 : _GEN_156; // @[FFT.scala 105:{12,12}]
  wire [16:0] _GEN_158 = 7'h1d == _wnList_T[6:0] ? _wnList_res_re_T_751 : _GEN_157; // @[FFT.scala 105:{12,12}]
  wire [16:0] _GEN_159 = 7'h1e == _wnList_T[6:0] ? _wnList_res_re_T_759 : _GEN_158; // @[FFT.scala 105:{12,12}]
  wire [16:0] _GEN_160 = 7'h1f == _wnList_T[6:0] ? _wnList_res_re_T_767 : _GEN_159; // @[FFT.scala 105:{12,12}]
  wire [16:0] _GEN_161 = 7'h20 == _wnList_T[6:0] ? _wnList_res_re_T_775 : _GEN_160; // @[FFT.scala 105:{12,12}]
  wire [16:0] _GEN_162 = 7'h21 == _wnList_T[6:0] ? _wnList_res_re_T_783 : _GEN_161; // @[FFT.scala 105:{12,12}]
  wire [16:0] _GEN_163 = 7'h22 == _wnList_T[6:0] ? _wnList_res_re_T_791 : _GEN_162; // @[FFT.scala 105:{12,12}]
  wire [16:0] _GEN_164 = 7'h23 == _wnList_T[6:0] ? _wnList_res_re_T_799 : _GEN_163; // @[FFT.scala 105:{12,12}]
  wire [16:0] _GEN_165 = 7'h24 == _wnList_T[6:0] ? _wnList_res_re_T_807 : _GEN_164; // @[FFT.scala 105:{12,12}]
  wire [16:0] _GEN_166 = 7'h25 == _wnList_T[6:0] ? _wnList_res_re_T_815 : _GEN_165; // @[FFT.scala 105:{12,12}]
  wire [16:0] _GEN_167 = 7'h26 == _wnList_T[6:0] ? _wnList_res_re_T_823 : _GEN_166; // @[FFT.scala 105:{12,12}]
  wire [16:0] _GEN_168 = 7'h27 == _wnList_T[6:0] ? _wnList_res_re_T_831 : _GEN_167; // @[FFT.scala 105:{12,12}]
  wire [16:0] _GEN_169 = 7'h28 == _wnList_T[6:0] ? _wnList_res_re_T_839 : _GEN_168; // @[FFT.scala 105:{12,12}]
  wire [16:0] _GEN_170 = 7'h29 == _wnList_T[6:0] ? _wnList_res_re_T_847 : _GEN_169; // @[FFT.scala 105:{12,12}]
  wire [16:0] _GEN_171 = 7'h2a == _wnList_T[6:0] ? _wnList_res_re_T_855 : _GEN_170; // @[FFT.scala 105:{12,12}]
  wire [16:0] _GEN_172 = 7'h2b == _wnList_T[6:0] ? _wnList_res_re_T_863 : _GEN_171; // @[FFT.scala 105:{12,12}]
  wire [16:0] _GEN_173 = 7'h2c == _wnList_T[6:0] ? _wnList_res_re_T_871 : _GEN_172; // @[FFT.scala 105:{12,12}]
  wire [16:0] _GEN_174 = 7'h2d == _wnList_T[6:0] ? _wnList_res_re_T_879 : _GEN_173; // @[FFT.scala 105:{12,12}]
  wire [16:0] _GEN_175 = 7'h2e == _wnList_T[6:0] ? _wnList_res_re_T_887 : _GEN_174; // @[FFT.scala 105:{12,12}]
  wire [16:0] _GEN_176 = 7'h2f == _wnList_T[6:0] ? _wnList_res_re_T_895 : _GEN_175; // @[FFT.scala 105:{12,12}]
  wire [16:0] _GEN_177 = 7'h30 == _wnList_T[6:0] ? _wnList_res_re_T_903 : _GEN_176; // @[FFT.scala 105:{12,12}]
  wire [16:0] _GEN_178 = 7'h31 == _wnList_T[6:0] ? _wnList_res_re_T_911 : _GEN_177; // @[FFT.scala 105:{12,12}]
  wire [16:0] _GEN_179 = 7'h32 == _wnList_T[6:0] ? _wnList_res_re_T_919 : _GEN_178; // @[FFT.scala 105:{12,12}]
  wire [16:0] _GEN_180 = 7'h33 == _wnList_T[6:0] ? _wnList_res_re_T_927 : _GEN_179; // @[FFT.scala 105:{12,12}]
  wire [16:0] _GEN_181 = 7'h34 == _wnList_T[6:0] ? _wnList_res_re_T_935 : _GEN_180; // @[FFT.scala 105:{12,12}]
  wire [16:0] _GEN_182 = 7'h35 == _wnList_T[6:0] ? _wnList_res_re_T_943 : _GEN_181; // @[FFT.scala 105:{12,12}]
  wire [16:0] _GEN_183 = 7'h36 == _wnList_T[6:0] ? _wnList_res_re_T_951 : _GEN_182; // @[FFT.scala 105:{12,12}]
  wire [16:0] _GEN_184 = 7'h37 == _wnList_T[6:0] ? _wnList_res_re_T_959 : _GEN_183; // @[FFT.scala 105:{12,12}]
  wire [16:0] _GEN_185 = 7'h38 == _wnList_T[6:0] ? _wnList_res_re_T_967 : _GEN_184; // @[FFT.scala 105:{12,12}]
  wire [16:0] _GEN_186 = 7'h39 == _wnList_T[6:0] ? _wnList_res_re_T_975 : _GEN_185; // @[FFT.scala 105:{12,12}]
  wire [16:0] _GEN_187 = 7'h3a == _wnList_T[6:0] ? _wnList_res_re_T_983 : _GEN_186; // @[FFT.scala 105:{12,12}]
  wire [16:0] _GEN_188 = 7'h3b == _wnList_T[6:0] ? _wnList_res_re_T_991 : _GEN_187; // @[FFT.scala 105:{12,12}]
  wire [16:0] _GEN_189 = 7'h3c == _wnList_T[6:0] ? _wnList_res_re_T_999 : _GEN_188; // @[FFT.scala 105:{12,12}]
  wire [16:0] _GEN_190 = 7'h3d == _wnList_T[6:0] ? _wnList_res_re_T_1007 : _GEN_189; // @[FFT.scala 105:{12,12}]
  wire [16:0] _GEN_191 = 7'h3e == _wnList_T[6:0] ? _wnList_res_re_T_1015 : _GEN_190; // @[FFT.scala 105:{12,12}]
  wire [16:0] _GEN_192 = 7'h3f == _wnList_T[6:0] ? _wnList_res_re_T_1023 : _GEN_191; // @[FFT.scala 105:{12,12}]
  wire [16:0] _GEN_193 = 7'h40 == _wnList_T[6:0] ? _wnList_res_im_T_519 : _GEN_192; // @[FFT.scala 105:{12,12}]
  wire [16:0] _GEN_194 = 7'h41 == _wnList_T[6:0] ? _wnList_res_re_T_1023 : _GEN_193; // @[FFT.scala 105:{12,12}]
  wire [16:0] _GEN_195 = 7'h42 == _wnList_T[6:0] ? _wnList_res_re_T_1015 : _GEN_194; // @[FFT.scala 105:{12,12}]
  wire [16:0] _GEN_196 = 7'h43 == _wnList_T[6:0] ? _wnList_res_re_T_1007 : _GEN_195; // @[FFT.scala 105:{12,12}]
  wire [16:0] _GEN_197 = 7'h44 == _wnList_T[6:0] ? _wnList_res_re_T_999 : _GEN_196; // @[FFT.scala 105:{12,12}]
  wire [16:0] _GEN_198 = 7'h45 == _wnList_T[6:0] ? _wnList_res_re_T_991 : _GEN_197; // @[FFT.scala 105:{12,12}]
  wire [16:0] _GEN_199 = 7'h46 == _wnList_T[6:0] ? _wnList_res_re_T_983 : _GEN_198; // @[FFT.scala 105:{12,12}]
  wire [16:0] _GEN_200 = 7'h47 == _wnList_T[6:0] ? _wnList_res_re_T_975 : _GEN_199; // @[FFT.scala 105:{12,12}]
  wire [16:0] _GEN_201 = 7'h48 == _wnList_T[6:0] ? _wnList_res_re_T_967 : _GEN_200; // @[FFT.scala 105:{12,12}]
  wire [16:0] _GEN_202 = 7'h49 == _wnList_T[6:0] ? _wnList_res_re_T_959 : _GEN_201; // @[FFT.scala 105:{12,12}]
  wire [16:0] _GEN_203 = 7'h4a == _wnList_T[6:0] ? _wnList_res_re_T_951 : _GEN_202; // @[FFT.scala 105:{12,12}]
  wire [16:0] _GEN_204 = 7'h4b == _wnList_T[6:0] ? _wnList_res_re_T_943 : _GEN_203; // @[FFT.scala 105:{12,12}]
  wire [16:0] _GEN_205 = 7'h4c == _wnList_T[6:0] ? _wnList_res_re_T_935 : _GEN_204; // @[FFT.scala 105:{12,12}]
  wire [16:0] _GEN_206 = 7'h4d == _wnList_T[6:0] ? _wnList_res_re_T_927 : _GEN_205; // @[FFT.scala 105:{12,12}]
  wire [16:0] _GEN_207 = 7'h4e == _wnList_T[6:0] ? _wnList_res_re_T_919 : _GEN_206; // @[FFT.scala 105:{12,12}]
  wire [16:0] _GEN_208 = 7'h4f == _wnList_T[6:0] ? _wnList_res_re_T_911 : _GEN_207; // @[FFT.scala 105:{12,12}]
  wire [16:0] _GEN_209 = 7'h50 == _wnList_T[6:0] ? _wnList_res_re_T_903 : _GEN_208; // @[FFT.scala 105:{12,12}]
  wire [16:0] _GEN_210 = 7'h51 == _wnList_T[6:0] ? _wnList_res_re_T_895 : _GEN_209; // @[FFT.scala 105:{12,12}]
  wire [16:0] _GEN_211 = 7'h52 == _wnList_T[6:0] ? _wnList_res_re_T_887 : _GEN_210; // @[FFT.scala 105:{12,12}]
  wire [16:0] _GEN_212 = 7'h53 == _wnList_T[6:0] ? _wnList_res_re_T_879 : _GEN_211; // @[FFT.scala 105:{12,12}]
  wire [16:0] _GEN_213 = 7'h54 == _wnList_T[6:0] ? _wnList_res_re_T_871 : _GEN_212; // @[FFT.scala 105:{12,12}]
  wire [16:0] _GEN_214 = 7'h55 == _wnList_T[6:0] ? _wnList_res_re_T_863 : _GEN_213; // @[FFT.scala 105:{12,12}]
  wire [16:0] _GEN_215 = 7'h56 == _wnList_T[6:0] ? _wnList_res_re_T_855 : _GEN_214; // @[FFT.scala 105:{12,12}]
  wire [16:0] _GEN_216 = 7'h57 == _wnList_T[6:0] ? _wnList_res_re_T_847 : _GEN_215; // @[FFT.scala 105:{12,12}]
  wire [16:0] _GEN_217 = 7'h58 == _wnList_T[6:0] ? _wnList_res_re_T_839 : _GEN_216; // @[FFT.scala 105:{12,12}]
  wire [16:0] _GEN_218 = 7'h59 == _wnList_T[6:0] ? _wnList_res_re_T_831 : _GEN_217; // @[FFT.scala 105:{12,12}]
  wire [16:0] _GEN_219 = 7'h5a == _wnList_T[6:0] ? _wnList_res_re_T_823 : _GEN_218; // @[FFT.scala 105:{12,12}]
  wire [16:0] _GEN_220 = 7'h5b == _wnList_T[6:0] ? _wnList_res_re_T_815 : _GEN_219; // @[FFT.scala 105:{12,12}]
  wire [16:0] _GEN_221 = 7'h5c == _wnList_T[6:0] ? _wnList_res_re_T_807 : _GEN_220; // @[FFT.scala 105:{12,12}]
  wire [16:0] _GEN_222 = 7'h5d == _wnList_T[6:0] ? _wnList_res_re_T_799 : _GEN_221; // @[FFT.scala 105:{12,12}]
  wire [16:0] _GEN_223 = 7'h5e == _wnList_T[6:0] ? _wnList_res_re_T_791 : _GEN_222; // @[FFT.scala 105:{12,12}]
  wire [16:0] _GEN_224 = 7'h5f == _wnList_T[6:0] ? _wnList_res_re_T_783 : _GEN_223; // @[FFT.scala 105:{12,12}]
  wire [16:0] _GEN_225 = 7'h60 == _wnList_T[6:0] ? _wnList_res_re_T_775 : _GEN_224; // @[FFT.scala 105:{12,12}]
  wire [16:0] _GEN_226 = 7'h61 == _wnList_T[6:0] ? _wnList_res_re_T_767 : _GEN_225; // @[FFT.scala 105:{12,12}]
  wire [16:0] _GEN_227 = 7'h62 == _wnList_T[6:0] ? _wnList_res_re_T_759 : _GEN_226; // @[FFT.scala 105:{12,12}]
  wire [16:0] _GEN_228 = 7'h63 == _wnList_T[6:0] ? _wnList_res_re_T_751 : _GEN_227; // @[FFT.scala 105:{12,12}]
  wire [16:0] _GEN_229 = 7'h64 == _wnList_T[6:0] ? _wnList_res_re_T_743 : _GEN_228; // @[FFT.scala 105:{12,12}]
  wire [16:0] _GEN_230 = 7'h65 == _wnList_T[6:0] ? _wnList_res_re_T_735 : _GEN_229; // @[FFT.scala 105:{12,12}]
  wire [16:0] _GEN_231 = 7'h66 == _wnList_T[6:0] ? _wnList_res_re_T_727 : _GEN_230; // @[FFT.scala 105:{12,12}]
  wire [16:0] _GEN_232 = 7'h67 == _wnList_T[6:0] ? _wnList_res_re_T_719 : _GEN_231; // @[FFT.scala 105:{12,12}]
  wire [16:0] _GEN_233 = 7'h68 == _wnList_T[6:0] ? _wnList_res_re_T_711 : _GEN_232; // @[FFT.scala 105:{12,12}]
  wire [16:0] _GEN_234 = 7'h69 == _wnList_T[6:0] ? _wnList_res_re_T_703 : _GEN_233; // @[FFT.scala 105:{12,12}]
  wire [16:0] _GEN_235 = 7'h6a == _wnList_T[6:0] ? _wnList_res_re_T_695 : _GEN_234; // @[FFT.scala 105:{12,12}]
  wire [16:0] _GEN_236 = 7'h6b == _wnList_T[6:0] ? _wnList_res_re_T_687 : _GEN_235; // @[FFT.scala 105:{12,12}]
  wire [16:0] _GEN_237 = 7'h6c == _wnList_T[6:0] ? _wnList_res_re_T_679 : _GEN_236; // @[FFT.scala 105:{12,12}]
  wire [16:0] _GEN_238 = 7'h6d == _wnList_T[6:0] ? _wnList_res_re_T_671 : _GEN_237; // @[FFT.scala 105:{12,12}]
  wire [16:0] _GEN_239 = 7'h6e == _wnList_T[6:0] ? _wnList_res_re_T_663 : _GEN_238; // @[FFT.scala 105:{12,12}]
  wire [16:0] _GEN_240 = 7'h6f == _wnList_T[6:0] ? _wnList_res_re_T_655 : _GEN_239; // @[FFT.scala 105:{12,12}]
  wire [16:0] _GEN_241 = 7'h70 == _wnList_T[6:0] ? _wnList_res_re_T_647 : _GEN_240; // @[FFT.scala 105:{12,12}]
  wire [16:0] _GEN_242 = 7'h71 == _wnList_T[6:0] ? _wnList_res_re_T_639 : _GEN_241; // @[FFT.scala 105:{12,12}]
  wire [16:0] _GEN_243 = 7'h72 == _wnList_T[6:0] ? _wnList_res_re_T_631 : _GEN_242; // @[FFT.scala 105:{12,12}]
  wire [16:0] _GEN_244 = 7'h73 == _wnList_T[6:0] ? _wnList_res_re_T_623 : _GEN_243; // @[FFT.scala 105:{12,12}]
  wire [16:0] _GEN_245 = 7'h74 == _wnList_T[6:0] ? _wnList_res_re_T_615 : _GEN_244; // @[FFT.scala 105:{12,12}]
  wire [16:0] _GEN_246 = 7'h75 == _wnList_T[6:0] ? _wnList_res_re_T_607 : _GEN_245; // @[FFT.scala 105:{12,12}]
  wire [16:0] _GEN_247 = 7'h76 == _wnList_T[6:0] ? _wnList_res_re_T_599 : _GEN_246; // @[FFT.scala 105:{12,12}]
  wire [16:0] _GEN_248 = 7'h77 == _wnList_T[6:0] ? _wnList_res_re_T_591 : _GEN_247; // @[FFT.scala 105:{12,12}]
  wire [16:0] _GEN_249 = 7'h78 == _wnList_T[6:0] ? _wnList_res_re_T_583 : _GEN_248; // @[FFT.scala 105:{12,12}]
  wire [16:0] _GEN_250 = 7'h79 == _wnList_T[6:0] ? _wnList_res_re_T_575 : _GEN_249; // @[FFT.scala 105:{12,12}]
  wire [16:0] _GEN_251 = 7'h7a == _wnList_T[6:0] ? _wnList_res_re_T_567 : _GEN_250; // @[FFT.scala 105:{12,12}]
  wire [16:0] _GEN_252 = 7'h7b == _wnList_T[6:0] ? _wnList_res_re_T_559 : _GEN_251; // @[FFT.scala 105:{12,12}]
  wire [16:0] _GEN_253 = 7'h7c == _wnList_T[6:0] ? _wnList_res_re_T_551 : _GEN_252; // @[FFT.scala 105:{12,12}]
  wire [16:0] _GEN_254 = 7'h7d == _wnList_T[6:0] ? _wnList_res_re_T_543 : _GEN_253; // @[FFT.scala 105:{12,12}]
  wire [16:0] _GEN_255 = 7'h7e == _wnList_T[6:0] ? _wnList_res_re_T_535 : _GEN_254; // @[FFT.scala 105:{12,12}]
  wire [5:0] wnCtrl_1 = cnt_0[5:0]; // @[FFT.scala 131:23]
  wire [6:0] _wnList_T_2 = {{1'd0}, wnCtrl_1}; // @[FFT.scala 135:96]
  wire [16:0] _GEN_258 = 6'h1 == _wnList_T_2[5:0] ? _wnList_res_re_T_23 : _wnList_res_re_T_7; // @[FFT.scala 104:{12,12}]
  wire [16:0] _GEN_259 = 6'h2 == _wnList_T_2[5:0] ? _wnList_res_re_T_39 : _GEN_258; // @[FFT.scala 104:{12,12}]
  wire [16:0] _GEN_260 = 6'h3 == _wnList_T_2[5:0] ? _wnList_res_re_T_55 : _GEN_259; // @[FFT.scala 104:{12,12}]
  wire [16:0] _GEN_261 = 6'h4 == _wnList_T_2[5:0] ? _wnList_res_re_T_71 : _GEN_260; // @[FFT.scala 104:{12,12}]
  wire [16:0] _GEN_262 = 6'h5 == _wnList_T_2[5:0] ? _wnList_res_re_T_87 : _GEN_261; // @[FFT.scala 104:{12,12}]
  wire [16:0] _GEN_263 = 6'h6 == _wnList_T_2[5:0] ? _wnList_res_re_T_103 : _GEN_262; // @[FFT.scala 104:{12,12}]
  wire [16:0] _GEN_264 = 6'h7 == _wnList_T_2[5:0] ? _wnList_res_re_T_119 : _GEN_263; // @[FFT.scala 104:{12,12}]
  wire [16:0] _GEN_265 = 6'h8 == _wnList_T_2[5:0] ? _wnList_res_re_T_135 : _GEN_264; // @[FFT.scala 104:{12,12}]
  wire [16:0] _GEN_266 = 6'h9 == _wnList_T_2[5:0] ? _wnList_res_re_T_151 : _GEN_265; // @[FFT.scala 104:{12,12}]
  wire [16:0] _GEN_267 = 6'ha == _wnList_T_2[5:0] ? _wnList_res_re_T_167 : _GEN_266; // @[FFT.scala 104:{12,12}]
  wire [16:0] _GEN_268 = 6'hb == _wnList_T_2[5:0] ? _wnList_res_re_T_183 : _GEN_267; // @[FFT.scala 104:{12,12}]
  wire [16:0] _GEN_269 = 6'hc == _wnList_T_2[5:0] ? _wnList_res_re_T_199 : _GEN_268; // @[FFT.scala 104:{12,12}]
  wire [16:0] _GEN_270 = 6'hd == _wnList_T_2[5:0] ? _wnList_res_re_T_215 : _GEN_269; // @[FFT.scala 104:{12,12}]
  wire [16:0] _GEN_271 = 6'he == _wnList_T_2[5:0] ? _wnList_res_re_T_231 : _GEN_270; // @[FFT.scala 104:{12,12}]
  wire [16:0] _GEN_272 = 6'hf == _wnList_T_2[5:0] ? _wnList_res_re_T_247 : _GEN_271; // @[FFT.scala 104:{12,12}]
  wire [16:0] _GEN_273 = 6'h10 == _wnList_T_2[5:0] ? _wnList_res_re_T_263 : _GEN_272; // @[FFT.scala 104:{12,12}]
  wire [16:0] _GEN_274 = 6'h11 == _wnList_T_2[5:0] ? _wnList_res_re_T_279 : _GEN_273; // @[FFT.scala 104:{12,12}]
  wire [16:0] _GEN_275 = 6'h12 == _wnList_T_2[5:0] ? _wnList_res_re_T_295 : _GEN_274; // @[FFT.scala 104:{12,12}]
  wire [16:0] _GEN_276 = 6'h13 == _wnList_T_2[5:0] ? _wnList_res_re_T_311 : _GEN_275; // @[FFT.scala 104:{12,12}]
  wire [16:0] _GEN_277 = 6'h14 == _wnList_T_2[5:0] ? _wnList_res_re_T_327 : _GEN_276; // @[FFT.scala 104:{12,12}]
  wire [16:0] _GEN_278 = 6'h15 == _wnList_T_2[5:0] ? _wnList_res_re_T_343 : _GEN_277; // @[FFT.scala 104:{12,12}]
  wire [16:0] _GEN_279 = 6'h16 == _wnList_T_2[5:0] ? _wnList_res_re_T_359 : _GEN_278; // @[FFT.scala 104:{12,12}]
  wire [16:0] _GEN_280 = 6'h17 == _wnList_T_2[5:0] ? _wnList_res_re_T_375 : _GEN_279; // @[FFT.scala 104:{12,12}]
  wire [16:0] _GEN_281 = 6'h18 == _wnList_T_2[5:0] ? _wnList_res_re_T_391 : _GEN_280; // @[FFT.scala 104:{12,12}]
  wire [16:0] _GEN_282 = 6'h19 == _wnList_T_2[5:0] ? _wnList_res_re_T_407 : _GEN_281; // @[FFT.scala 104:{12,12}]
  wire [16:0] _GEN_283 = 6'h1a == _wnList_T_2[5:0] ? _wnList_res_re_T_423 : _GEN_282; // @[FFT.scala 104:{12,12}]
  wire [16:0] _GEN_284 = 6'h1b == _wnList_T_2[5:0] ? _wnList_res_re_T_439 : _GEN_283; // @[FFT.scala 104:{12,12}]
  wire [16:0] _GEN_285 = 6'h1c == _wnList_T_2[5:0] ? _wnList_res_re_T_455 : _GEN_284; // @[FFT.scala 104:{12,12}]
  wire [16:0] _GEN_286 = 6'h1d == _wnList_T_2[5:0] ? _wnList_res_re_T_471 : _GEN_285; // @[FFT.scala 104:{12,12}]
  wire [16:0] _GEN_287 = 6'h1e == _wnList_T_2[5:0] ? _wnList_res_re_T_487 : _GEN_286; // @[FFT.scala 104:{12,12}]
  wire [16:0] _GEN_288 = 6'h1f == _wnList_T_2[5:0] ? _wnList_res_re_T_503 : _GEN_287; // @[FFT.scala 104:{12,12}]
  wire [16:0] _GEN_289 = 6'h20 == _wnList_T_2[5:0] ? _wnList_res_re_T_519 : _GEN_288; // @[FFT.scala 104:{12,12}]
  wire [16:0] _GEN_290 = 6'h21 == _wnList_T_2[5:0] ? _wnList_res_re_T_535 : _GEN_289; // @[FFT.scala 104:{12,12}]
  wire [16:0] _GEN_291 = 6'h22 == _wnList_T_2[5:0] ? _wnList_res_re_T_551 : _GEN_290; // @[FFT.scala 104:{12,12}]
  wire [16:0] _GEN_292 = 6'h23 == _wnList_T_2[5:0] ? _wnList_res_re_T_567 : _GEN_291; // @[FFT.scala 104:{12,12}]
  wire [16:0] _GEN_293 = 6'h24 == _wnList_T_2[5:0] ? _wnList_res_re_T_583 : _GEN_292; // @[FFT.scala 104:{12,12}]
  wire [16:0] _GEN_294 = 6'h25 == _wnList_T_2[5:0] ? _wnList_res_re_T_599 : _GEN_293; // @[FFT.scala 104:{12,12}]
  wire [16:0] _GEN_295 = 6'h26 == _wnList_T_2[5:0] ? _wnList_res_re_T_615 : _GEN_294; // @[FFT.scala 104:{12,12}]
  wire [16:0] _GEN_296 = 6'h27 == _wnList_T_2[5:0] ? _wnList_res_re_T_631 : _GEN_295; // @[FFT.scala 104:{12,12}]
  wire [16:0] _GEN_297 = 6'h28 == _wnList_T_2[5:0] ? _wnList_res_re_T_647 : _GEN_296; // @[FFT.scala 104:{12,12}]
  wire [16:0] _GEN_298 = 6'h29 == _wnList_T_2[5:0] ? _wnList_res_re_T_663 : _GEN_297; // @[FFT.scala 104:{12,12}]
  wire [16:0] _GEN_299 = 6'h2a == _wnList_T_2[5:0] ? _wnList_res_re_T_679 : _GEN_298; // @[FFT.scala 104:{12,12}]
  wire [16:0] _GEN_300 = 6'h2b == _wnList_T_2[5:0] ? _wnList_res_re_T_695 : _GEN_299; // @[FFT.scala 104:{12,12}]
  wire [16:0] _GEN_301 = 6'h2c == _wnList_T_2[5:0] ? _wnList_res_re_T_711 : _GEN_300; // @[FFT.scala 104:{12,12}]
  wire [16:0] _GEN_302 = 6'h2d == _wnList_T_2[5:0] ? _wnList_res_re_T_727 : _GEN_301; // @[FFT.scala 104:{12,12}]
  wire [16:0] _GEN_303 = 6'h2e == _wnList_T_2[5:0] ? _wnList_res_re_T_743 : _GEN_302; // @[FFT.scala 104:{12,12}]
  wire [16:0] _GEN_304 = 6'h2f == _wnList_T_2[5:0] ? _wnList_res_re_T_759 : _GEN_303; // @[FFT.scala 104:{12,12}]
  wire [16:0] _GEN_305 = 6'h30 == _wnList_T_2[5:0] ? _wnList_res_re_T_775 : _GEN_304; // @[FFT.scala 104:{12,12}]
  wire [16:0] _GEN_306 = 6'h31 == _wnList_T_2[5:0] ? _wnList_res_re_T_791 : _GEN_305; // @[FFT.scala 104:{12,12}]
  wire [16:0] _GEN_307 = 6'h32 == _wnList_T_2[5:0] ? _wnList_res_re_T_807 : _GEN_306; // @[FFT.scala 104:{12,12}]
  wire [16:0] _GEN_308 = 6'h33 == _wnList_T_2[5:0] ? _wnList_res_re_T_823 : _GEN_307; // @[FFT.scala 104:{12,12}]
  wire [16:0] _GEN_309 = 6'h34 == _wnList_T_2[5:0] ? _wnList_res_re_T_839 : _GEN_308; // @[FFT.scala 104:{12,12}]
  wire [16:0] _GEN_310 = 6'h35 == _wnList_T_2[5:0] ? _wnList_res_re_T_855 : _GEN_309; // @[FFT.scala 104:{12,12}]
  wire [16:0] _GEN_311 = 6'h36 == _wnList_T_2[5:0] ? _wnList_res_re_T_871 : _GEN_310; // @[FFT.scala 104:{12,12}]
  wire [16:0] _GEN_312 = 6'h37 == _wnList_T_2[5:0] ? _wnList_res_re_T_887 : _GEN_311; // @[FFT.scala 104:{12,12}]
  wire [16:0] _GEN_313 = 6'h38 == _wnList_T_2[5:0] ? _wnList_res_re_T_903 : _GEN_312; // @[FFT.scala 104:{12,12}]
  wire [16:0] _GEN_314 = 6'h39 == _wnList_T_2[5:0] ? _wnList_res_re_T_919 : _GEN_313; // @[FFT.scala 104:{12,12}]
  wire [16:0] _GEN_315 = 6'h3a == _wnList_T_2[5:0] ? _wnList_res_re_T_935 : _GEN_314; // @[FFT.scala 104:{12,12}]
  wire [16:0] _GEN_316 = 6'h3b == _wnList_T_2[5:0] ? _wnList_res_re_T_951 : _GEN_315; // @[FFT.scala 104:{12,12}]
  wire [16:0] _GEN_317 = 6'h3c == _wnList_T_2[5:0] ? _wnList_res_re_T_967 : _GEN_316; // @[FFT.scala 104:{12,12}]
  wire [16:0] _GEN_318 = 6'h3d == _wnList_T_2[5:0] ? _wnList_res_re_T_983 : _GEN_317; // @[FFT.scala 104:{12,12}]
  wire [16:0] _GEN_319 = 6'h3e == _wnList_T_2[5:0] ? _wnList_res_re_T_999 : _GEN_318; // @[FFT.scala 104:{12,12}]
  wire [16:0] _GEN_322 = 6'h1 == _wnList_T_2[5:0] ? _wnList_res_re_T_535 : _wnList_res_re_T_519; // @[FFT.scala 105:{12,12}]
  wire [16:0] _GEN_323 = 6'h2 == _wnList_T_2[5:0] ? _wnList_res_re_T_551 : _GEN_322; // @[FFT.scala 105:{12,12}]
  wire [16:0] _GEN_324 = 6'h3 == _wnList_T_2[5:0] ? _wnList_res_re_T_567 : _GEN_323; // @[FFT.scala 105:{12,12}]
  wire [16:0] _GEN_325 = 6'h4 == _wnList_T_2[5:0] ? _wnList_res_re_T_583 : _GEN_324; // @[FFT.scala 105:{12,12}]
  wire [16:0] _GEN_326 = 6'h5 == _wnList_T_2[5:0] ? _wnList_res_re_T_599 : _GEN_325; // @[FFT.scala 105:{12,12}]
  wire [16:0] _GEN_327 = 6'h6 == _wnList_T_2[5:0] ? _wnList_res_re_T_615 : _GEN_326; // @[FFT.scala 105:{12,12}]
  wire [16:0] _GEN_328 = 6'h7 == _wnList_T_2[5:0] ? _wnList_res_re_T_631 : _GEN_327; // @[FFT.scala 105:{12,12}]
  wire [16:0] _GEN_329 = 6'h8 == _wnList_T_2[5:0] ? _wnList_res_re_T_647 : _GEN_328; // @[FFT.scala 105:{12,12}]
  wire [16:0] _GEN_330 = 6'h9 == _wnList_T_2[5:0] ? _wnList_res_re_T_663 : _GEN_329; // @[FFT.scala 105:{12,12}]
  wire [16:0] _GEN_331 = 6'ha == _wnList_T_2[5:0] ? _wnList_res_re_T_679 : _GEN_330; // @[FFT.scala 105:{12,12}]
  wire [16:0] _GEN_332 = 6'hb == _wnList_T_2[5:0] ? _wnList_res_re_T_695 : _GEN_331; // @[FFT.scala 105:{12,12}]
  wire [16:0] _GEN_333 = 6'hc == _wnList_T_2[5:0] ? _wnList_res_re_T_711 : _GEN_332; // @[FFT.scala 105:{12,12}]
  wire [16:0] _GEN_334 = 6'hd == _wnList_T_2[5:0] ? _wnList_res_re_T_727 : _GEN_333; // @[FFT.scala 105:{12,12}]
  wire [16:0] _GEN_335 = 6'he == _wnList_T_2[5:0] ? _wnList_res_re_T_743 : _GEN_334; // @[FFT.scala 105:{12,12}]
  wire [16:0] _GEN_336 = 6'hf == _wnList_T_2[5:0] ? _wnList_res_re_T_759 : _GEN_335; // @[FFT.scala 105:{12,12}]
  wire [16:0] _GEN_337 = 6'h10 == _wnList_T_2[5:0] ? _wnList_res_re_T_775 : _GEN_336; // @[FFT.scala 105:{12,12}]
  wire [16:0] _GEN_338 = 6'h11 == _wnList_T_2[5:0] ? _wnList_res_re_T_791 : _GEN_337; // @[FFT.scala 105:{12,12}]
  wire [16:0] _GEN_339 = 6'h12 == _wnList_T_2[5:0] ? _wnList_res_re_T_807 : _GEN_338; // @[FFT.scala 105:{12,12}]
  wire [16:0] _GEN_340 = 6'h13 == _wnList_T_2[5:0] ? _wnList_res_re_T_823 : _GEN_339; // @[FFT.scala 105:{12,12}]
  wire [16:0] _GEN_341 = 6'h14 == _wnList_T_2[5:0] ? _wnList_res_re_T_839 : _GEN_340; // @[FFT.scala 105:{12,12}]
  wire [16:0] _GEN_342 = 6'h15 == _wnList_T_2[5:0] ? _wnList_res_re_T_855 : _GEN_341; // @[FFT.scala 105:{12,12}]
  wire [16:0] _GEN_343 = 6'h16 == _wnList_T_2[5:0] ? _wnList_res_re_T_871 : _GEN_342; // @[FFT.scala 105:{12,12}]
  wire [16:0] _GEN_344 = 6'h17 == _wnList_T_2[5:0] ? _wnList_res_re_T_887 : _GEN_343; // @[FFT.scala 105:{12,12}]
  wire [16:0] _GEN_345 = 6'h18 == _wnList_T_2[5:0] ? _wnList_res_re_T_903 : _GEN_344; // @[FFT.scala 105:{12,12}]
  wire [16:0] _GEN_346 = 6'h19 == _wnList_T_2[5:0] ? _wnList_res_re_T_919 : _GEN_345; // @[FFT.scala 105:{12,12}]
  wire [16:0] _GEN_347 = 6'h1a == _wnList_T_2[5:0] ? _wnList_res_re_T_935 : _GEN_346; // @[FFT.scala 105:{12,12}]
  wire [16:0] _GEN_348 = 6'h1b == _wnList_T_2[5:0] ? _wnList_res_re_T_951 : _GEN_347; // @[FFT.scala 105:{12,12}]
  wire [16:0] _GEN_349 = 6'h1c == _wnList_T_2[5:0] ? _wnList_res_re_T_967 : _GEN_348; // @[FFT.scala 105:{12,12}]
  wire [16:0] _GEN_350 = 6'h1d == _wnList_T_2[5:0] ? _wnList_res_re_T_983 : _GEN_349; // @[FFT.scala 105:{12,12}]
  wire [16:0] _GEN_351 = 6'h1e == _wnList_T_2[5:0] ? _wnList_res_re_T_999 : _GEN_350; // @[FFT.scala 105:{12,12}]
  wire [16:0] _GEN_352 = 6'h1f == _wnList_T_2[5:0] ? _wnList_res_re_T_1015 : _GEN_351; // @[FFT.scala 105:{12,12}]
  wire [16:0] _GEN_353 = 6'h20 == _wnList_T_2[5:0] ? _wnList_res_im_T_519 : _GEN_352; // @[FFT.scala 105:{12,12}]
  wire [16:0] _GEN_354 = 6'h21 == _wnList_T_2[5:0] ? _wnList_res_re_T_1015 : _GEN_353; // @[FFT.scala 105:{12,12}]
  wire [16:0] _GEN_355 = 6'h22 == _wnList_T_2[5:0] ? _wnList_res_re_T_999 : _GEN_354; // @[FFT.scala 105:{12,12}]
  wire [16:0] _GEN_356 = 6'h23 == _wnList_T_2[5:0] ? _wnList_res_re_T_983 : _GEN_355; // @[FFT.scala 105:{12,12}]
  wire [16:0] _GEN_357 = 6'h24 == _wnList_T_2[5:0] ? _wnList_res_re_T_967 : _GEN_356; // @[FFT.scala 105:{12,12}]
  wire [16:0] _GEN_358 = 6'h25 == _wnList_T_2[5:0] ? _wnList_res_re_T_951 : _GEN_357; // @[FFT.scala 105:{12,12}]
  wire [16:0] _GEN_359 = 6'h26 == _wnList_T_2[5:0] ? _wnList_res_re_T_935 : _GEN_358; // @[FFT.scala 105:{12,12}]
  wire [16:0] _GEN_360 = 6'h27 == _wnList_T_2[5:0] ? _wnList_res_re_T_919 : _GEN_359; // @[FFT.scala 105:{12,12}]
  wire [16:0] _GEN_361 = 6'h28 == _wnList_T_2[5:0] ? _wnList_res_re_T_903 : _GEN_360; // @[FFT.scala 105:{12,12}]
  wire [16:0] _GEN_362 = 6'h29 == _wnList_T_2[5:0] ? _wnList_res_re_T_887 : _GEN_361; // @[FFT.scala 105:{12,12}]
  wire [16:0] _GEN_363 = 6'h2a == _wnList_T_2[5:0] ? _wnList_res_re_T_871 : _GEN_362; // @[FFT.scala 105:{12,12}]
  wire [16:0] _GEN_364 = 6'h2b == _wnList_T_2[5:0] ? _wnList_res_re_T_855 : _GEN_363; // @[FFT.scala 105:{12,12}]
  wire [16:0] _GEN_365 = 6'h2c == _wnList_T_2[5:0] ? _wnList_res_re_T_839 : _GEN_364; // @[FFT.scala 105:{12,12}]
  wire [16:0] _GEN_366 = 6'h2d == _wnList_T_2[5:0] ? _wnList_res_re_T_823 : _GEN_365; // @[FFT.scala 105:{12,12}]
  wire [16:0] _GEN_367 = 6'h2e == _wnList_T_2[5:0] ? _wnList_res_re_T_807 : _GEN_366; // @[FFT.scala 105:{12,12}]
  wire [16:0] _GEN_368 = 6'h2f == _wnList_T_2[5:0] ? _wnList_res_re_T_791 : _GEN_367; // @[FFT.scala 105:{12,12}]
  wire [16:0] _GEN_369 = 6'h30 == _wnList_T_2[5:0] ? _wnList_res_re_T_775 : _GEN_368; // @[FFT.scala 105:{12,12}]
  wire [16:0] _GEN_370 = 6'h31 == _wnList_T_2[5:0] ? _wnList_res_re_T_759 : _GEN_369; // @[FFT.scala 105:{12,12}]
  wire [16:0] _GEN_371 = 6'h32 == _wnList_T_2[5:0] ? _wnList_res_re_T_743 : _GEN_370; // @[FFT.scala 105:{12,12}]
  wire [16:0] _GEN_372 = 6'h33 == _wnList_T_2[5:0] ? _wnList_res_re_T_727 : _GEN_371; // @[FFT.scala 105:{12,12}]
  wire [16:0] _GEN_373 = 6'h34 == _wnList_T_2[5:0] ? _wnList_res_re_T_711 : _GEN_372; // @[FFT.scala 105:{12,12}]
  wire [16:0] _GEN_374 = 6'h35 == _wnList_T_2[5:0] ? _wnList_res_re_T_695 : _GEN_373; // @[FFT.scala 105:{12,12}]
  wire [16:0] _GEN_375 = 6'h36 == _wnList_T_2[5:0] ? _wnList_res_re_T_679 : _GEN_374; // @[FFT.scala 105:{12,12}]
  wire [16:0] _GEN_376 = 6'h37 == _wnList_T_2[5:0] ? _wnList_res_re_T_663 : _GEN_375; // @[FFT.scala 105:{12,12}]
  wire [16:0] _GEN_377 = 6'h38 == _wnList_T_2[5:0] ? _wnList_res_re_T_647 : _GEN_376; // @[FFT.scala 105:{12,12}]
  wire [16:0] _GEN_378 = 6'h39 == _wnList_T_2[5:0] ? _wnList_res_re_T_631 : _GEN_377; // @[FFT.scala 105:{12,12}]
  wire [16:0] _GEN_379 = 6'h3a == _wnList_T_2[5:0] ? _wnList_res_re_T_615 : _GEN_378; // @[FFT.scala 105:{12,12}]
  wire [16:0] _GEN_380 = 6'h3b == _wnList_T_2[5:0] ? _wnList_res_re_T_599 : _GEN_379; // @[FFT.scala 105:{12,12}]
  wire [16:0] _GEN_381 = 6'h3c == _wnList_T_2[5:0] ? _wnList_res_re_T_583 : _GEN_380; // @[FFT.scala 105:{12,12}]
  wire [16:0] _GEN_382 = 6'h3d == _wnList_T_2[5:0] ? _wnList_res_re_T_567 : _GEN_381; // @[FFT.scala 105:{12,12}]
  wire [16:0] _GEN_383 = 6'h3e == _wnList_T_2[5:0] ? _wnList_res_re_T_551 : _GEN_382; // @[FFT.scala 105:{12,12}]
  wire [4:0] wnCtrl_2 = cnt_0[4:0]; // @[FFT.scala 131:23]
  wire [5:0] _wnList_T_4 = {{1'd0}, wnCtrl_2}; // @[FFT.scala 135:96]
  wire [16:0] _GEN_386 = 5'h1 == _wnList_T_4[4:0] ? _wnList_res_re_T_39 : _wnList_res_re_T_7; // @[FFT.scala 104:{12,12}]
  wire [16:0] _GEN_387 = 5'h2 == _wnList_T_4[4:0] ? _wnList_res_re_T_71 : _GEN_386; // @[FFT.scala 104:{12,12}]
  wire [16:0] _GEN_388 = 5'h3 == _wnList_T_4[4:0] ? _wnList_res_re_T_103 : _GEN_387; // @[FFT.scala 104:{12,12}]
  wire [16:0] _GEN_389 = 5'h4 == _wnList_T_4[4:0] ? _wnList_res_re_T_135 : _GEN_388; // @[FFT.scala 104:{12,12}]
  wire [16:0] _GEN_390 = 5'h5 == _wnList_T_4[4:0] ? _wnList_res_re_T_167 : _GEN_389; // @[FFT.scala 104:{12,12}]
  wire [16:0] _GEN_391 = 5'h6 == _wnList_T_4[4:0] ? _wnList_res_re_T_199 : _GEN_390; // @[FFT.scala 104:{12,12}]
  wire [16:0] _GEN_392 = 5'h7 == _wnList_T_4[4:0] ? _wnList_res_re_T_231 : _GEN_391; // @[FFT.scala 104:{12,12}]
  wire [16:0] _GEN_393 = 5'h8 == _wnList_T_4[4:0] ? _wnList_res_re_T_263 : _GEN_392; // @[FFT.scala 104:{12,12}]
  wire [16:0] _GEN_394 = 5'h9 == _wnList_T_4[4:0] ? _wnList_res_re_T_295 : _GEN_393; // @[FFT.scala 104:{12,12}]
  wire [16:0] _GEN_395 = 5'ha == _wnList_T_4[4:0] ? _wnList_res_re_T_327 : _GEN_394; // @[FFT.scala 104:{12,12}]
  wire [16:0] _GEN_396 = 5'hb == _wnList_T_4[4:0] ? _wnList_res_re_T_359 : _GEN_395; // @[FFT.scala 104:{12,12}]
  wire [16:0] _GEN_397 = 5'hc == _wnList_T_4[4:0] ? _wnList_res_re_T_391 : _GEN_396; // @[FFT.scala 104:{12,12}]
  wire [16:0] _GEN_398 = 5'hd == _wnList_T_4[4:0] ? _wnList_res_re_T_423 : _GEN_397; // @[FFT.scala 104:{12,12}]
  wire [16:0] _GEN_399 = 5'he == _wnList_T_4[4:0] ? _wnList_res_re_T_455 : _GEN_398; // @[FFT.scala 104:{12,12}]
  wire [16:0] _GEN_400 = 5'hf == _wnList_T_4[4:0] ? _wnList_res_re_T_487 : _GEN_399; // @[FFT.scala 104:{12,12}]
  wire [16:0] _GEN_401 = 5'h10 == _wnList_T_4[4:0] ? _wnList_res_re_T_519 : _GEN_400; // @[FFT.scala 104:{12,12}]
  wire [16:0] _GEN_402 = 5'h11 == _wnList_T_4[4:0] ? _wnList_res_re_T_551 : _GEN_401; // @[FFT.scala 104:{12,12}]
  wire [16:0] _GEN_403 = 5'h12 == _wnList_T_4[4:0] ? _wnList_res_re_T_583 : _GEN_402; // @[FFT.scala 104:{12,12}]
  wire [16:0] _GEN_404 = 5'h13 == _wnList_T_4[4:0] ? _wnList_res_re_T_615 : _GEN_403; // @[FFT.scala 104:{12,12}]
  wire [16:0] _GEN_405 = 5'h14 == _wnList_T_4[4:0] ? _wnList_res_re_T_647 : _GEN_404; // @[FFT.scala 104:{12,12}]
  wire [16:0] _GEN_406 = 5'h15 == _wnList_T_4[4:0] ? _wnList_res_re_T_679 : _GEN_405; // @[FFT.scala 104:{12,12}]
  wire [16:0] _GEN_407 = 5'h16 == _wnList_T_4[4:0] ? _wnList_res_re_T_711 : _GEN_406; // @[FFT.scala 104:{12,12}]
  wire [16:0] _GEN_408 = 5'h17 == _wnList_T_4[4:0] ? _wnList_res_re_T_743 : _GEN_407; // @[FFT.scala 104:{12,12}]
  wire [16:0] _GEN_409 = 5'h18 == _wnList_T_4[4:0] ? _wnList_res_re_T_775 : _GEN_408; // @[FFT.scala 104:{12,12}]
  wire [16:0] _GEN_410 = 5'h19 == _wnList_T_4[4:0] ? _wnList_res_re_T_807 : _GEN_409; // @[FFT.scala 104:{12,12}]
  wire [16:0] _GEN_411 = 5'h1a == _wnList_T_4[4:0] ? _wnList_res_re_T_839 : _GEN_410; // @[FFT.scala 104:{12,12}]
  wire [16:0] _GEN_412 = 5'h1b == _wnList_T_4[4:0] ? _wnList_res_re_T_871 : _GEN_411; // @[FFT.scala 104:{12,12}]
  wire [16:0] _GEN_413 = 5'h1c == _wnList_T_4[4:0] ? _wnList_res_re_T_903 : _GEN_412; // @[FFT.scala 104:{12,12}]
  wire [16:0] _GEN_414 = 5'h1d == _wnList_T_4[4:0] ? _wnList_res_re_T_935 : _GEN_413; // @[FFT.scala 104:{12,12}]
  wire [16:0] _GEN_415 = 5'h1e == _wnList_T_4[4:0] ? _wnList_res_re_T_967 : _GEN_414; // @[FFT.scala 104:{12,12}]
  wire [16:0] _GEN_418 = 5'h1 == _wnList_T_4[4:0] ? _wnList_res_re_T_551 : _wnList_res_re_T_519; // @[FFT.scala 105:{12,12}]
  wire [16:0] _GEN_419 = 5'h2 == _wnList_T_4[4:0] ? _wnList_res_re_T_583 : _GEN_418; // @[FFT.scala 105:{12,12}]
  wire [16:0] _GEN_420 = 5'h3 == _wnList_T_4[4:0] ? _wnList_res_re_T_615 : _GEN_419; // @[FFT.scala 105:{12,12}]
  wire [16:0] _GEN_421 = 5'h4 == _wnList_T_4[4:0] ? _wnList_res_re_T_647 : _GEN_420; // @[FFT.scala 105:{12,12}]
  wire [16:0] _GEN_422 = 5'h5 == _wnList_T_4[4:0] ? _wnList_res_re_T_679 : _GEN_421; // @[FFT.scala 105:{12,12}]
  wire [16:0] _GEN_423 = 5'h6 == _wnList_T_4[4:0] ? _wnList_res_re_T_711 : _GEN_422; // @[FFT.scala 105:{12,12}]
  wire [16:0] _GEN_424 = 5'h7 == _wnList_T_4[4:0] ? _wnList_res_re_T_743 : _GEN_423; // @[FFT.scala 105:{12,12}]
  wire [16:0] _GEN_425 = 5'h8 == _wnList_T_4[4:0] ? _wnList_res_re_T_775 : _GEN_424; // @[FFT.scala 105:{12,12}]
  wire [16:0] _GEN_426 = 5'h9 == _wnList_T_4[4:0] ? _wnList_res_re_T_807 : _GEN_425; // @[FFT.scala 105:{12,12}]
  wire [16:0] _GEN_427 = 5'ha == _wnList_T_4[4:0] ? _wnList_res_re_T_839 : _GEN_426; // @[FFT.scala 105:{12,12}]
  wire [16:0] _GEN_428 = 5'hb == _wnList_T_4[4:0] ? _wnList_res_re_T_871 : _GEN_427; // @[FFT.scala 105:{12,12}]
  wire [16:0] _GEN_429 = 5'hc == _wnList_T_4[4:0] ? _wnList_res_re_T_903 : _GEN_428; // @[FFT.scala 105:{12,12}]
  wire [16:0] _GEN_430 = 5'hd == _wnList_T_4[4:0] ? _wnList_res_re_T_935 : _GEN_429; // @[FFT.scala 105:{12,12}]
  wire [16:0] _GEN_431 = 5'he == _wnList_T_4[4:0] ? _wnList_res_re_T_967 : _GEN_430; // @[FFT.scala 105:{12,12}]
  wire [16:0] _GEN_432 = 5'hf == _wnList_T_4[4:0] ? _wnList_res_re_T_999 : _GEN_431; // @[FFT.scala 105:{12,12}]
  wire [16:0] _GEN_433 = 5'h10 == _wnList_T_4[4:0] ? _wnList_res_im_T_519 : _GEN_432; // @[FFT.scala 105:{12,12}]
  wire [16:0] _GEN_434 = 5'h11 == _wnList_T_4[4:0] ? _wnList_res_re_T_999 : _GEN_433; // @[FFT.scala 105:{12,12}]
  wire [16:0] _GEN_435 = 5'h12 == _wnList_T_4[4:0] ? _wnList_res_re_T_967 : _GEN_434; // @[FFT.scala 105:{12,12}]
  wire [16:0] _GEN_436 = 5'h13 == _wnList_T_4[4:0] ? _wnList_res_re_T_935 : _GEN_435; // @[FFT.scala 105:{12,12}]
  wire [16:0] _GEN_437 = 5'h14 == _wnList_T_4[4:0] ? _wnList_res_re_T_903 : _GEN_436; // @[FFT.scala 105:{12,12}]
  wire [16:0] _GEN_438 = 5'h15 == _wnList_T_4[4:0] ? _wnList_res_re_T_871 : _GEN_437; // @[FFT.scala 105:{12,12}]
  wire [16:0] _GEN_439 = 5'h16 == _wnList_T_4[4:0] ? _wnList_res_re_T_839 : _GEN_438; // @[FFT.scala 105:{12,12}]
  wire [16:0] _GEN_440 = 5'h17 == _wnList_T_4[4:0] ? _wnList_res_re_T_807 : _GEN_439; // @[FFT.scala 105:{12,12}]
  wire [16:0] _GEN_441 = 5'h18 == _wnList_T_4[4:0] ? _wnList_res_re_T_775 : _GEN_440; // @[FFT.scala 105:{12,12}]
  wire [16:0] _GEN_442 = 5'h19 == _wnList_T_4[4:0] ? _wnList_res_re_T_743 : _GEN_441; // @[FFT.scala 105:{12,12}]
  wire [16:0] _GEN_443 = 5'h1a == _wnList_T_4[4:0] ? _wnList_res_re_T_711 : _GEN_442; // @[FFT.scala 105:{12,12}]
  wire [16:0] _GEN_444 = 5'h1b == _wnList_T_4[4:0] ? _wnList_res_re_T_679 : _GEN_443; // @[FFT.scala 105:{12,12}]
  wire [16:0] _GEN_445 = 5'h1c == _wnList_T_4[4:0] ? _wnList_res_re_T_647 : _GEN_444; // @[FFT.scala 105:{12,12}]
  wire [16:0] _GEN_446 = 5'h1d == _wnList_T_4[4:0] ? _wnList_res_re_T_615 : _GEN_445; // @[FFT.scala 105:{12,12}]
  wire [16:0] _GEN_447 = 5'h1e == _wnList_T_4[4:0] ? _wnList_res_re_T_583 : _GEN_446; // @[FFT.scala 105:{12,12}]
  wire [3:0] wnCtrl_3 = cnt_0[3:0]; // @[FFT.scala 131:23]
  wire [4:0] _wnList_T_6 = {{1'd0}, wnCtrl_3}; // @[FFT.scala 135:96]
  wire [16:0] _GEN_450 = 4'h1 == _wnList_T_6[3:0] ? _wnList_res_re_T_71 : _wnList_res_re_T_7; // @[FFT.scala 104:{12,12}]
  wire [16:0] _GEN_451 = 4'h2 == _wnList_T_6[3:0] ? _wnList_res_re_T_135 : _GEN_450; // @[FFT.scala 104:{12,12}]
  wire [16:0] _GEN_452 = 4'h3 == _wnList_T_6[3:0] ? _wnList_res_re_T_199 : _GEN_451; // @[FFT.scala 104:{12,12}]
  wire [16:0] _GEN_453 = 4'h4 == _wnList_T_6[3:0] ? _wnList_res_re_T_263 : _GEN_452; // @[FFT.scala 104:{12,12}]
  wire [16:0] _GEN_454 = 4'h5 == _wnList_T_6[3:0] ? _wnList_res_re_T_327 : _GEN_453; // @[FFT.scala 104:{12,12}]
  wire [16:0] _GEN_455 = 4'h6 == _wnList_T_6[3:0] ? _wnList_res_re_T_391 : _GEN_454; // @[FFT.scala 104:{12,12}]
  wire [16:0] _GEN_456 = 4'h7 == _wnList_T_6[3:0] ? _wnList_res_re_T_455 : _GEN_455; // @[FFT.scala 104:{12,12}]
  wire [16:0] _GEN_457 = 4'h8 == _wnList_T_6[3:0] ? _wnList_res_re_T_519 : _GEN_456; // @[FFT.scala 104:{12,12}]
  wire [16:0] _GEN_458 = 4'h9 == _wnList_T_6[3:0] ? _wnList_res_re_T_583 : _GEN_457; // @[FFT.scala 104:{12,12}]
  wire [16:0] _GEN_459 = 4'ha == _wnList_T_6[3:0] ? _wnList_res_re_T_647 : _GEN_458; // @[FFT.scala 104:{12,12}]
  wire [16:0] _GEN_460 = 4'hb == _wnList_T_6[3:0] ? _wnList_res_re_T_711 : _GEN_459; // @[FFT.scala 104:{12,12}]
  wire [16:0] _GEN_461 = 4'hc == _wnList_T_6[3:0] ? _wnList_res_re_T_775 : _GEN_460; // @[FFT.scala 104:{12,12}]
  wire [16:0] _GEN_462 = 4'hd == _wnList_T_6[3:0] ? _wnList_res_re_T_839 : _GEN_461; // @[FFT.scala 104:{12,12}]
  wire [16:0] _GEN_463 = 4'he == _wnList_T_6[3:0] ? _wnList_res_re_T_903 : _GEN_462; // @[FFT.scala 104:{12,12}]
  wire [16:0] _GEN_466 = 4'h1 == _wnList_T_6[3:0] ? _wnList_res_re_T_583 : _wnList_res_re_T_519; // @[FFT.scala 105:{12,12}]
  wire [16:0] _GEN_467 = 4'h2 == _wnList_T_6[3:0] ? _wnList_res_re_T_647 : _GEN_466; // @[FFT.scala 105:{12,12}]
  wire [16:0] _GEN_468 = 4'h3 == _wnList_T_6[3:0] ? _wnList_res_re_T_711 : _GEN_467; // @[FFT.scala 105:{12,12}]
  wire [16:0] _GEN_469 = 4'h4 == _wnList_T_6[3:0] ? _wnList_res_re_T_775 : _GEN_468; // @[FFT.scala 105:{12,12}]
  wire [16:0] _GEN_470 = 4'h5 == _wnList_T_6[3:0] ? _wnList_res_re_T_839 : _GEN_469; // @[FFT.scala 105:{12,12}]
  wire [16:0] _GEN_471 = 4'h6 == _wnList_T_6[3:0] ? _wnList_res_re_T_903 : _GEN_470; // @[FFT.scala 105:{12,12}]
  wire [16:0] _GEN_472 = 4'h7 == _wnList_T_6[3:0] ? _wnList_res_re_T_967 : _GEN_471; // @[FFT.scala 105:{12,12}]
  wire [16:0] _GEN_473 = 4'h8 == _wnList_T_6[3:0] ? _wnList_res_im_T_519 : _GEN_472; // @[FFT.scala 105:{12,12}]
  wire [16:0] _GEN_474 = 4'h9 == _wnList_T_6[3:0] ? _wnList_res_re_T_967 : _GEN_473; // @[FFT.scala 105:{12,12}]
  wire [16:0] _GEN_475 = 4'ha == _wnList_T_6[3:0] ? _wnList_res_re_T_903 : _GEN_474; // @[FFT.scala 105:{12,12}]
  wire [16:0] _GEN_476 = 4'hb == _wnList_T_6[3:0] ? _wnList_res_re_T_839 : _GEN_475; // @[FFT.scala 105:{12,12}]
  wire [16:0] _GEN_477 = 4'hc == _wnList_T_6[3:0] ? _wnList_res_re_T_775 : _GEN_476; // @[FFT.scala 105:{12,12}]
  wire [16:0] _GEN_478 = 4'hd == _wnList_T_6[3:0] ? _wnList_res_re_T_711 : _GEN_477; // @[FFT.scala 105:{12,12}]
  wire [16:0] _GEN_479 = 4'he == _wnList_T_6[3:0] ? _wnList_res_re_T_647 : _GEN_478; // @[FFT.scala 105:{12,12}]
  wire [2:0] wnCtrl_4 = cnt_0[2:0]; // @[FFT.scala 131:23]
  wire [3:0] _wnList_T_8 = {{1'd0}, wnCtrl_4}; // @[FFT.scala 135:96]
  wire [16:0] _GEN_482 = 3'h1 == _wnList_T_8[2:0] ? _wnList_res_re_T_135 : _wnList_res_re_T_7; // @[FFT.scala 104:{12,12}]
  wire [16:0] _GEN_483 = 3'h2 == _wnList_T_8[2:0] ? _wnList_res_re_T_263 : _GEN_482; // @[FFT.scala 104:{12,12}]
  wire [16:0] _GEN_484 = 3'h3 == _wnList_T_8[2:0] ? _wnList_res_re_T_391 : _GEN_483; // @[FFT.scala 104:{12,12}]
  wire [16:0] _GEN_485 = 3'h4 == _wnList_T_8[2:0] ? _wnList_res_re_T_519 : _GEN_484; // @[FFT.scala 104:{12,12}]
  wire [16:0] _GEN_486 = 3'h5 == _wnList_T_8[2:0] ? _wnList_res_re_T_647 : _GEN_485; // @[FFT.scala 104:{12,12}]
  wire [16:0] _GEN_487 = 3'h6 == _wnList_T_8[2:0] ? _wnList_res_re_T_775 : _GEN_486; // @[FFT.scala 104:{12,12}]
  wire [16:0] _GEN_490 = 3'h1 == _wnList_T_8[2:0] ? _wnList_res_re_T_647 : _wnList_res_re_T_519; // @[FFT.scala 105:{12,12}]
  wire [16:0] _GEN_491 = 3'h2 == _wnList_T_8[2:0] ? _wnList_res_re_T_775 : _GEN_490; // @[FFT.scala 105:{12,12}]
  wire [16:0] _GEN_492 = 3'h3 == _wnList_T_8[2:0] ? _wnList_res_re_T_903 : _GEN_491; // @[FFT.scala 105:{12,12}]
  wire [16:0] _GEN_493 = 3'h4 == _wnList_T_8[2:0] ? _wnList_res_im_T_519 : _GEN_492; // @[FFT.scala 105:{12,12}]
  wire [16:0] _GEN_494 = 3'h5 == _wnList_T_8[2:0] ? _wnList_res_re_T_903 : _GEN_493; // @[FFT.scala 105:{12,12}]
  wire [16:0] _GEN_495 = 3'h6 == _wnList_T_8[2:0] ? _wnList_res_re_T_775 : _GEN_494; // @[FFT.scala 105:{12,12}]
  wire [1:0] wnCtrl_5 = cnt_0[1:0]; // @[FFT.scala 131:23]
  wire [2:0] _wnList_T_10 = {{1'd0}, wnCtrl_5}; // @[FFT.scala 135:96]
  wire [16:0] _GEN_498 = 2'h1 == _wnList_T_10[1:0] ? _wnList_res_re_T_263 : _wnList_res_re_T_7; // @[FFT.scala 104:{12,12}]
  wire [16:0] _GEN_499 = 2'h2 == _wnList_T_10[1:0] ? _wnList_res_re_T_519 : _GEN_498; // @[FFT.scala 104:{12,12}]
  wire [16:0] _GEN_502 = 2'h1 == _wnList_T_10[1:0] ? _wnList_res_re_T_775 : _wnList_res_re_T_519; // @[FFT.scala 105:{12,12}]
  wire [16:0] _GEN_503 = 2'h2 == _wnList_T_10[1:0] ? _wnList_res_im_T_519 : _GEN_502; // @[FFT.scala 105:{12,12}]
  wire  wnCtrl_6 = cnt_0[0]; // @[FFT.scala 131:23]
  wire [1:0] _wnList_T_12 = {{1'd0}, wnCtrl_6}; // @[FFT.scala 135:96]
  wire [31:0] _T_1 = {io_dIn_0_re,io_dIn_0_im}; // @[FFT.scala 170:91]
  wire [31:0] _T_4 = {io_dIn_1_re,io_dIn_1_im}; // @[FFT.scala 170:91]
  reg [8:0] io_dout_valid_REG; // @[FFT.scala 179:27]
  wire [16:0] datao_0_re = dataotemp_inst_io_out_0_re; // @[FFT.scala 124:22 141:9]
  wire [16:0] datao_0_im = dataotemp_inst_io_out_0_im; // @[FFT.scala 124:22 141:9]
  wire [33:0] _T_7 = {datao_0_re,datao_0_im}; // @[FFT.scala 181:96]
  reg [15:0] REG_re; // @[FFT.scala 181:64]
  reg [15:0] REG_im; // @[FFT.scala 181:64]
  wire [16:0] datao_1_re = dataotemp_inst_io_out_1_re; // @[FFT.scala 124:22 141:9]
  wire [16:0] datao_1_im = dataotemp_inst_io_out_1_im; // @[FFT.scala 124:22 141:9]
  wire [33:0] _T_10 = {datao_1_re,datao_1_im}; // @[FFT.scala 181:96]
  reg [15:0] REG_1_re; // @[FFT.scala 181:64]
  reg [15:0] REG_1_im; // @[FFT.scala 181:64]
  ButterflyMul inst ( // @[Modules.scala 287:22]
    .io_in_0_re(inst_io_in_0_re),
    .io_in_0_im(inst_io_in_0_im),
    .io_in_1_re(inst_io_in_1_re),
    .io_in_1_im(inst_io_in_1_im),
    .io_out_0_re(inst_io_out_0_re),
    .io_out_0_im(inst_io_out_0_im),
    .io_out_1_re(inst_io_out_1_re),
    .io_out_1_im(inst_io_out_1_im),
    .io_wn_0_re(inst_io_wn_0_re),
    .io_wn_0_im(inst_io_wn_0_im)
  );
  ButterflyMul inst_1 ( // @[Modules.scala 287:22]
    .io_in_0_re(inst_1_io_in_0_re),
    .io_in_0_im(inst_1_io_in_0_im),
    .io_in_1_re(inst_1_io_in_1_re),
    .io_in_1_im(inst_1_io_in_1_im),
    .io_out_0_re(inst_1_io_out_0_re),
    .io_out_0_im(inst_1_io_out_0_im),
    .io_out_1_re(inst_1_io_out_1_re),
    .io_out_1_im(inst_1_io_out_1_im),
    .io_wn_0_re(inst_1_io_wn_0_re),
    .io_wn_0_im(inst_1_io_wn_0_im)
  );
  ButterflyMul inst_2 ( // @[Modules.scala 287:22]
    .io_in_0_re(inst_2_io_in_0_re),
    .io_in_0_im(inst_2_io_in_0_im),
    .io_in_1_re(inst_2_io_in_1_re),
    .io_in_1_im(inst_2_io_in_1_im),
    .io_out_0_re(inst_2_io_out_0_re),
    .io_out_0_im(inst_2_io_out_0_im),
    .io_out_1_re(inst_2_io_out_1_re),
    .io_out_1_im(inst_2_io_out_1_im),
    .io_wn_0_re(inst_2_io_wn_0_re),
    .io_wn_0_im(inst_2_io_wn_0_im)
  );
  ButterflyMul inst_3 ( // @[Modules.scala 287:22]
    .io_in_0_re(inst_3_io_in_0_re),
    .io_in_0_im(inst_3_io_in_0_im),
    .io_in_1_re(inst_3_io_in_1_re),
    .io_in_1_im(inst_3_io_in_1_im),
    .io_out_0_re(inst_3_io_out_0_re),
    .io_out_0_im(inst_3_io_out_0_im),
    .io_out_1_re(inst_3_io_out_1_re),
    .io_out_1_im(inst_3_io_out_1_im),
    .io_wn_0_re(inst_3_io_wn_0_re),
    .io_wn_0_im(inst_3_io_wn_0_im)
  );
  ButterflyMul inst_4 ( // @[Modules.scala 287:22]
    .io_in_0_re(inst_4_io_in_0_re),
    .io_in_0_im(inst_4_io_in_0_im),
    .io_in_1_re(inst_4_io_in_1_re),
    .io_in_1_im(inst_4_io_in_1_im),
    .io_out_0_re(inst_4_io_out_0_re),
    .io_out_0_im(inst_4_io_out_0_im),
    .io_out_1_re(inst_4_io_out_1_re),
    .io_out_1_im(inst_4_io_out_1_im),
    .io_wn_0_re(inst_4_io_wn_0_re),
    .io_wn_0_im(inst_4_io_wn_0_im)
  );
  ButterflyMul inst_5 ( // @[Modules.scala 287:22]
    .io_in_0_re(inst_5_io_in_0_re),
    .io_in_0_im(inst_5_io_in_0_im),
    .io_in_1_re(inst_5_io_in_1_re),
    .io_in_1_im(inst_5_io_in_1_im),
    .io_out_0_re(inst_5_io_out_0_re),
    .io_out_0_im(inst_5_io_out_0_im),
    .io_out_1_re(inst_5_io_out_1_re),
    .io_out_1_im(inst_5_io_out_1_im),
    .io_wn_0_re(inst_5_io_wn_0_re),
    .io_wn_0_im(inst_5_io_wn_0_im)
  );
  ButterflyMul inst_6 ( // @[Modules.scala 287:22]
    .io_in_0_re(inst_6_io_in_0_re),
    .io_in_0_im(inst_6_io_in_0_im),
    .io_in_1_re(inst_6_io_in_1_re),
    .io_in_1_im(inst_6_io_in_1_im),
    .io_out_0_re(inst_6_io_out_0_re),
    .io_out_0_im(inst_6_io_out_0_im),
    .io_out_1_re(inst_6_io_out_1_re),
    .io_out_1_im(inst_6_io_out_1_im),
    .io_wn_0_re(inst_6_io_wn_0_re),
    .io_wn_0_im(inst_6_io_wn_0_im)
  );
  ButterflyAdd dataotemp_inst ( // @[Modules.scala 213:22]
    .io_in_0_re(dataotemp_inst_io_in_0_re),
    .io_in_0_im(dataotemp_inst_io_in_0_im),
    .io_in_1_re(dataotemp_inst_io_in_1_re),
    .io_in_1_im(dataotemp_inst_io_in_1_im),
    .io_out_0_re(dataotemp_inst_io_out_0_re),
    .io_out_0_im(dataotemp_inst_io_out_0_im),
    .io_out_1_re(dataotemp_inst_io_out_1_re),
    .io_out_1_im(dataotemp_inst_io_out_1_im)
  );
  Switch inst_7 ( // @[Modules.scala 311:22]
    .clock(inst_7_clock),
    .io_in_0_re(inst_7_io_in_0_re),
    .io_in_0_im(inst_7_io_in_0_im),
    .io_in_1_re(inst_7_io_in_1_re),
    .io_in_1_im(inst_7_io_in_1_im),
    .io_out_0_re(inst_7_io_out_0_re),
    .io_out_0_im(inst_7_io_out_0_im),
    .io_out_1_re(inst_7_io_out_1_re),
    .io_out_1_im(inst_7_io_out_1_im),
    .io_sel(inst_7_io_sel)
  );
  Switch_1 inst_8 ( // @[Modules.scala 311:22]
    .clock(inst_8_clock),
    .io_in_0_re(inst_8_io_in_0_re),
    .io_in_0_im(inst_8_io_in_0_im),
    .io_in_1_re(inst_8_io_in_1_re),
    .io_in_1_im(inst_8_io_in_1_im),
    .io_out_0_re(inst_8_io_out_0_re),
    .io_out_0_im(inst_8_io_out_0_im),
    .io_out_1_re(inst_8_io_out_1_re),
    .io_out_1_im(inst_8_io_out_1_im),
    .io_sel(inst_8_io_sel)
  );
  Switch_2 inst_9 ( // @[Modules.scala 311:22]
    .clock(inst_9_clock),
    .io_in_0_re(inst_9_io_in_0_re),
    .io_in_0_im(inst_9_io_in_0_im),
    .io_in_1_re(inst_9_io_in_1_re),
    .io_in_1_im(inst_9_io_in_1_im),
    .io_out_0_re(inst_9_io_out_0_re),
    .io_out_0_im(inst_9_io_out_0_im),
    .io_out_1_re(inst_9_io_out_1_re),
    .io_out_1_im(inst_9_io_out_1_im),
    .io_sel(inst_9_io_sel)
  );
  Switch_3 inst_10 ( // @[Modules.scala 311:22]
    .clock(inst_10_clock),
    .io_in_0_re(inst_10_io_in_0_re),
    .io_in_0_im(inst_10_io_in_0_im),
    .io_in_1_re(inst_10_io_in_1_re),
    .io_in_1_im(inst_10_io_in_1_im),
    .io_out_0_re(inst_10_io_out_0_re),
    .io_out_0_im(inst_10_io_out_0_im),
    .io_out_1_re(inst_10_io_out_1_re),
    .io_out_1_im(inst_10_io_out_1_im),
    .io_sel(inst_10_io_sel)
  );
  Switch_4 inst_11 ( // @[Modules.scala 311:22]
    .clock(inst_11_clock),
    .io_in_0_re(inst_11_io_in_0_re),
    .io_in_0_im(inst_11_io_in_0_im),
    .io_in_1_re(inst_11_io_in_1_re),
    .io_in_1_im(inst_11_io_in_1_im),
    .io_out_0_re(inst_11_io_out_0_re),
    .io_out_0_im(inst_11_io_out_0_im),
    .io_out_1_re(inst_11_io_out_1_re),
    .io_out_1_im(inst_11_io_out_1_im),
    .io_sel(inst_11_io_sel)
  );
  Switch_5 inst_12 ( // @[Modules.scala 311:22]
    .clock(inst_12_clock),
    .io_in_0_re(inst_12_io_in_0_re),
    .io_in_0_im(inst_12_io_in_0_im),
    .io_in_1_re(inst_12_io_in_1_re),
    .io_in_1_im(inst_12_io_in_1_im),
    .io_out_0_re(inst_12_io_out_0_re),
    .io_out_0_im(inst_12_io_out_0_im),
    .io_out_1_re(inst_12_io_out_1_re),
    .io_out_1_im(inst_12_io_out_1_im),
    .io_sel(inst_12_io_sel)
  );
  Switch_6 inst_13 ( // @[Modules.scala 311:22]
    .clock(inst_13_clock),
    .io_in_0_re(inst_13_io_in_0_re),
    .io_in_0_im(inst_13_io_in_0_im),
    .io_in_1_re(inst_13_io_in_1_re),
    .io_in_1_im(inst_13_io_in_1_im),
    .io_out_0_re(inst_13_io_out_0_re),
    .io_out_0_im(inst_13_io_out_0_im),
    .io_out_1_re(inst_13_io_out_1_re),
    .io_out_1_im(inst_13_io_out_1_im),
    .io_sel(inst_13_io_sel)
  );
  ComplexRecode inst_14 ( // @[Modules.scala 40:22]
    .io_in_re(inst_14_io_in_re),
    .io_in_im(inst_14_io_in_im),
    .io_out_re(inst_14_io_out_re),
    .io_out_im(inst_14_io_out_im)
  );
  ComplexRecode inst_15 ( // @[Modules.scala 40:22]
    .io_in_re(inst_15_io_in_re),
    .io_in_im(inst_15_io_in_im),
    .io_out_re(inst_15_io_out_re),
    .io_out_im(inst_15_io_out_im)
  );
  ComplexDecode inst_16 ( // @[Modules.scala 56:22]
    .io_in_re(inst_16_io_in_re),
    .io_in_im(inst_16_io_in_im),
    .io_out_re(inst_16_io_out_re),
    .io_out_im(inst_16_io_out_im)
  );
  ComplexDecode inst_17 ( // @[Modules.scala 56:22]
    .io_in_re(inst_17_io_in_re),
    .io_in_im(inst_17_io_in_im),
    .io_out_re(inst_17_io_out_re),
    .io_out_im(inst_17_io_out_im)
  );
  assign io_dOut_0_re = REG_re; // @[FFT.scala 181:13]
  assign io_dOut_0_im = REG_im; // @[FFT.scala 181:13]
  assign io_dOut_1_re = REG_1_re; // @[FFT.scala 181:13]
  assign io_dOut_1_im = REG_1_im; // @[FFT.scala 181:13]
  assign io_dout_valid = io_dout_valid_REG == 9'h7f; // @[FFT.scala 179:36]
  assign io_busy = cnt_0 != 9'h0; // @[FFT.scala 114:21]
  assign inst_io_in_0_re = inst_14_io_out_re; // @[FFT.scala 122:65 170:19]
  assign inst_io_in_0_im = inst_14_io_out_im; // @[FFT.scala 122:65 170:19]
  assign inst_io_in_1_re = inst_15_io_out_re; // @[FFT.scala 122:65 170:19]
  assign inst_io_in_1_im = inst_15_io_out_im; // @[FFT.scala 122:65 170:19]
  assign inst_io_wn_0_re = 7'h7f == _wnList_T[6:0] ? _wnList_res_re_T_1023 : _GEN_127; // @[FFT.scala 104:{12,12}]
  assign inst_io_wn_0_im = 7'h7f == _wnList_T[6:0] ? _wnList_res_re_T_527 : _GEN_255; // @[FFT.scala 105:{12,12}]
  assign inst_1_io_in_0_re = inst_7_io_out_0_re; // @[FFT.scala 122:65 164:54]
  assign inst_1_io_in_0_im = inst_7_io_out_0_im; // @[FFT.scala 122:65 164:54]
  assign inst_1_io_in_1_re = inst_7_io_out_1_re; // @[FFT.scala 122:65 164:54]
  assign inst_1_io_in_1_im = inst_7_io_out_1_im; // @[FFT.scala 122:65 164:54]
  assign inst_1_io_wn_0_re = 6'h3f == _wnList_T_2[5:0] ? _wnList_res_re_T_1015 : _GEN_319; // @[FFT.scala 104:{12,12}]
  assign inst_1_io_wn_0_im = 6'h3f == _wnList_T_2[5:0] ? _wnList_res_re_T_535 : _GEN_383; // @[FFT.scala 105:{12,12}]
  assign inst_2_io_in_0_re = inst_8_io_out_0_re; // @[FFT.scala 122:65 164:54]
  assign inst_2_io_in_0_im = inst_8_io_out_0_im; // @[FFT.scala 122:65 164:54]
  assign inst_2_io_in_1_re = inst_8_io_out_1_re; // @[FFT.scala 122:65 164:54]
  assign inst_2_io_in_1_im = inst_8_io_out_1_im; // @[FFT.scala 122:65 164:54]
  assign inst_2_io_wn_0_re = 5'h1f == _wnList_T_4[4:0] ? _wnList_res_re_T_999 : _GEN_415; // @[FFT.scala 104:{12,12}]
  assign inst_2_io_wn_0_im = 5'h1f == _wnList_T_4[4:0] ? _wnList_res_re_T_551 : _GEN_447; // @[FFT.scala 105:{12,12}]
  assign inst_3_io_in_0_re = inst_9_io_out_0_re; // @[FFT.scala 122:65 164:54]
  assign inst_3_io_in_0_im = inst_9_io_out_0_im; // @[FFT.scala 122:65 164:54]
  assign inst_3_io_in_1_re = inst_9_io_out_1_re; // @[FFT.scala 122:65 164:54]
  assign inst_3_io_in_1_im = inst_9_io_out_1_im; // @[FFT.scala 122:65 164:54]
  assign inst_3_io_wn_0_re = 4'hf == _wnList_T_6[3:0] ? _wnList_res_re_T_967 : _GEN_463; // @[FFT.scala 104:{12,12}]
  assign inst_3_io_wn_0_im = 4'hf == _wnList_T_6[3:0] ? _wnList_res_re_T_583 : _GEN_479; // @[FFT.scala 105:{12,12}]
  assign inst_4_io_in_0_re = inst_10_io_out_0_re; // @[FFT.scala 122:65 164:54]
  assign inst_4_io_in_0_im = inst_10_io_out_0_im; // @[FFT.scala 122:65 164:54]
  assign inst_4_io_in_1_re = inst_10_io_out_1_re; // @[FFT.scala 122:65 164:54]
  assign inst_4_io_in_1_im = inst_10_io_out_1_im; // @[FFT.scala 122:65 164:54]
  assign inst_4_io_wn_0_re = 3'h7 == _wnList_T_8[2:0] ? _wnList_res_re_T_903 : _GEN_487; // @[FFT.scala 104:{12,12}]
  assign inst_4_io_wn_0_im = 3'h7 == _wnList_T_8[2:0] ? _wnList_res_re_T_647 : _GEN_495; // @[FFT.scala 105:{12,12}]
  assign inst_5_io_in_0_re = inst_11_io_out_0_re; // @[FFT.scala 122:65 164:54]
  assign inst_5_io_in_0_im = inst_11_io_out_0_im; // @[FFT.scala 122:65 164:54]
  assign inst_5_io_in_1_re = inst_11_io_out_1_re; // @[FFT.scala 122:65 164:54]
  assign inst_5_io_in_1_im = inst_11_io_out_1_im; // @[FFT.scala 122:65 164:54]
  assign inst_5_io_wn_0_re = 2'h3 == _wnList_T_10[1:0] ? _wnList_res_re_T_775 : _GEN_499; // @[FFT.scala 104:{12,12}]
  assign inst_5_io_wn_0_im = 2'h3 == _wnList_T_10[1:0] ? _wnList_res_re_T_775 : _GEN_503; // @[FFT.scala 105:{12,12}]
  assign inst_6_io_in_0_re = inst_12_io_out_0_re; // @[FFT.scala 122:65 164:54]
  assign inst_6_io_in_0_im = inst_12_io_out_0_im; // @[FFT.scala 122:65 164:54]
  assign inst_6_io_in_1_re = inst_12_io_out_1_re; // @[FFT.scala 122:65 164:54]
  assign inst_6_io_in_1_im = inst_12_io_out_1_im; // @[FFT.scala 122:65 164:54]
  assign inst_6_io_wn_0_re = _wnList_T_12[0] ? _wnList_res_re_T_519 : _wnList_res_re_T_7; // @[FFT.scala 104:{12,12}]
  assign inst_6_io_wn_0_im = _wnList_T_12[0] ? _wnList_res_im_T_519 : _wnList_res_re_T_519; // @[FFT.scala 105:{12,12}]
  assign dataotemp_inst_io_in_0_re = inst_13_io_out_0_re; // @[FFT.scala 122:65 164:54]
  assign dataotemp_inst_io_in_0_im = inst_13_io_out_0_im; // @[FFT.scala 122:65 164:54]
  assign dataotemp_inst_io_in_1_re = inst_13_io_out_1_re; // @[FFT.scala 122:65 164:54]
  assign dataotemp_inst_io_in_1_im = inst_13_io_out_1_im; // @[FFT.scala 122:65 164:54]
  assign inst_7_clock = clock;
  assign inst_7_io_in_0_re = inst_io_out_0_re; // @[FFT.scala 123:69 136:19]
  assign inst_7_io_in_0_im = inst_io_out_0_im; // @[FFT.scala 123:69 136:19]
  assign inst_7_io_in_1_re = inst_io_out_1_re; // @[FFT.scala 123:69 136:19]
  assign inst_7_io_in_1_im = inst_io_out_1_im; // @[FFT.scala 123:69 136:19]
  assign inst_7_io_sel = cnt_0[6]; // @[FFT.scala 163:31]
  assign inst_8_clock = clock;
  assign inst_8_io_in_0_re = inst_1_io_out_0_re; // @[FFT.scala 123:69 136:19]
  assign inst_8_io_in_0_im = inst_1_io_out_0_im; // @[FFT.scala 123:69 136:19]
  assign inst_8_io_in_1_re = inst_1_io_out_1_re; // @[FFT.scala 123:69 136:19]
  assign inst_8_io_in_1_im = inst_1_io_out_1_im; // @[FFT.scala 123:69 136:19]
  assign inst_8_io_sel = cnt_0[5]; // @[FFT.scala 163:31]
  assign inst_9_clock = clock;
  assign inst_9_io_in_0_re = inst_2_io_out_0_re; // @[FFT.scala 123:69 136:19]
  assign inst_9_io_in_0_im = inst_2_io_out_0_im; // @[FFT.scala 123:69 136:19]
  assign inst_9_io_in_1_re = inst_2_io_out_1_re; // @[FFT.scala 123:69 136:19]
  assign inst_9_io_in_1_im = inst_2_io_out_1_im; // @[FFT.scala 123:69 136:19]
  assign inst_9_io_sel = cnt_0[4]; // @[FFT.scala 163:31]
  assign inst_10_clock = clock;
  assign inst_10_io_in_0_re = inst_3_io_out_0_re; // @[FFT.scala 123:69 136:19]
  assign inst_10_io_in_0_im = inst_3_io_out_0_im; // @[FFT.scala 123:69 136:19]
  assign inst_10_io_in_1_re = inst_3_io_out_1_re; // @[FFT.scala 123:69 136:19]
  assign inst_10_io_in_1_im = inst_3_io_out_1_im; // @[FFT.scala 123:69 136:19]
  assign inst_10_io_sel = cnt_0[3]; // @[FFT.scala 163:31]
  assign inst_11_clock = clock;
  assign inst_11_io_in_0_re = inst_4_io_out_0_re; // @[FFT.scala 123:69 136:19]
  assign inst_11_io_in_0_im = inst_4_io_out_0_im; // @[FFT.scala 123:69 136:19]
  assign inst_11_io_in_1_re = inst_4_io_out_1_re; // @[FFT.scala 123:69 136:19]
  assign inst_11_io_in_1_im = inst_4_io_out_1_im; // @[FFT.scala 123:69 136:19]
  assign inst_11_io_sel = cnt_0[2]; // @[FFT.scala 163:31]
  assign inst_12_clock = clock;
  assign inst_12_io_in_0_re = inst_5_io_out_0_re; // @[FFT.scala 123:69 136:19]
  assign inst_12_io_in_0_im = inst_5_io_out_0_im; // @[FFT.scala 123:69 136:19]
  assign inst_12_io_in_1_re = inst_5_io_out_1_re; // @[FFT.scala 123:69 136:19]
  assign inst_12_io_in_1_im = inst_5_io_out_1_im; // @[FFT.scala 123:69 136:19]
  assign inst_12_io_sel = cnt_0[1]; // @[FFT.scala 163:31]
  assign inst_13_clock = clock;
  assign inst_13_io_in_0_re = inst_6_io_out_0_re; // @[FFT.scala 123:69 136:19]
  assign inst_13_io_in_0_im = inst_6_io_out_0_im; // @[FFT.scala 123:69 136:19]
  assign inst_13_io_in_1_re = inst_6_io_out_1_re; // @[FFT.scala 123:69 136:19]
  assign inst_13_io_in_1_im = inst_6_io_out_1_im; // @[FFT.scala 123:69 136:19]
  assign inst_13_io_sel = cnt_0[0]; // @[FFT.scala 163:31]
  assign inst_14_io_in_re = _T_1[31:16]; // @[FFT.scala 170:91]
  assign inst_14_io_in_im = _T_1[15:0]; // @[FFT.scala 170:91]
  assign inst_15_io_in_re = _T_4[31:16]; // @[FFT.scala 170:91]
  assign inst_15_io_in_im = _T_4[15:0]; // @[FFT.scala 170:91]
  assign inst_16_io_in_re = _T_7[33:17]; // @[FFT.scala 181:96]
  assign inst_16_io_in_im = _T_7[16:0]; // @[FFT.scala 181:96]
  assign inst_17_io_in_re = _T_10[33:17]; // @[FFT.scala 181:96]
  assign inst_17_io_in_im = _T_10[16:0]; // @[FFT.scala 181:96]
  always @(posedge clock) begin
    if (reset) begin // @[FFT.scala 110:46]
      cnt_0 <= 9'h0; // @[FFT.scala 110:46]
    end else if (io_din_valid | busy) begin // @[FFT.scala 115:30]
      if (cnt_0 == 9'hff) begin // @[FFT.scala 116:18]
        cnt_0 <= 9'h0;
      end else begin
        cnt_0 <= _cnt_0_T_2;
      end
    end
    io_dout_valid_REG <= cnt_0; // @[FFT.scala 179:27]
    REG_re <= inst_16_io_out_re; // @[FFT.scala 181:64]
    REG_im <= inst_16_io_out_im; // @[FFT.scala 181:64]
    REG_1_re <= inst_17_io_out_re; // @[FFT.scala 181:64]
    REG_1_im <= inst_17_io_out_im; // @[FFT.scala 181:64]
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  cnt_0 = _RAND_0[8:0];
  _RAND_1 = {1{`RANDOM}};
  io_dout_valid_REG = _RAND_1[8:0];
  _RAND_2 = {1{`RANDOM}};
  REG_re = _RAND_2[15:0];
  _RAND_3 = {1{`RANDOM}};
  REG_im = _RAND_3[15:0];
  _RAND_4 = {1{`RANDOM}};
  REG_1_re = _RAND_4[15:0];
  _RAND_5 = {1{`RANDOM}};
  REG_1_im = _RAND_5[15:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module FFTtop(
  input         clock,
  input         reset,
  input  [15:0] io_dIn_0_re,
  input  [15:0] io_dIn_0_im,
  input  [15:0] io_dIn_1_re,
  input  [15:0] io_dIn_1_im,
  output [15:0] io_dOut_0_re,
  output [15:0] io_dOut_0_im,
  output [15:0] io_dOut_1_re,
  output [15:0] io_dOut_1_im,
  input         io_din_valid,
  output        io_dout_valid,
  output        io_busy
);
  wire  fft_clock; // @[Top.scala 15:19]
  wire  fft_reset; // @[Top.scala 15:19]
  wire [15:0] fft_io_dIn_0_re; // @[Top.scala 15:19]
  wire [15:0] fft_io_dIn_0_im; // @[Top.scala 15:19]
  wire [15:0] fft_io_dIn_1_re; // @[Top.scala 15:19]
  wire [15:0] fft_io_dIn_1_im; // @[Top.scala 15:19]
  wire [15:0] fft_io_dOut_0_re; // @[Top.scala 15:19]
  wire [15:0] fft_io_dOut_0_im; // @[Top.scala 15:19]
  wire [15:0] fft_io_dOut_1_re; // @[Top.scala 15:19]
  wire [15:0] fft_io_dOut_1_im; // @[Top.scala 15:19]
  wire  fft_io_din_valid; // @[Top.scala 15:19]
  wire  fft_io_dout_valid; // @[Top.scala 15:19]
  wire  fft_io_busy; // @[Top.scala 15:19]
  FFT fft ( // @[Top.scala 15:19]
    .clock(fft_clock),
    .reset(fft_reset),
    .io_dIn_0_re(fft_io_dIn_0_re),
    .io_dIn_0_im(fft_io_dIn_0_im),
    .io_dIn_1_re(fft_io_dIn_1_re),
    .io_dIn_1_im(fft_io_dIn_1_im),
    .io_dOut_0_re(fft_io_dOut_0_re),
    .io_dOut_0_im(fft_io_dOut_0_im),
    .io_dOut_1_re(fft_io_dOut_1_re),
    .io_dOut_1_im(fft_io_dOut_1_im),
    .io_din_valid(fft_io_din_valid),
    .io_dout_valid(fft_io_dout_valid),
    .io_busy(fft_io_busy)
  );
  assign io_dOut_0_re = fft_io_dOut_0_re; // @[Top.scala 27:13]
  assign io_dOut_0_im = fft_io_dOut_0_im; // @[Top.scala 27:13]
  assign io_dOut_1_re = fft_io_dOut_1_re; // @[Top.scala 27:13]
  assign io_dOut_1_im = fft_io_dOut_1_im; // @[Top.scala 27:13]
  assign io_dout_valid = fft_io_dout_valid; // @[Top.scala 28:19]
  assign io_busy = fft_io_busy; // @[Top.scala 29:13]
  assign fft_clock = clock;
  assign fft_reset = reset;
  assign fft_io_dIn_0_re = io_dIn_0_re; // @[Top.scala 16:14]
  assign fft_io_dIn_0_im = io_dIn_0_im; // @[Top.scala 16:14]
  assign fft_io_dIn_1_re = io_dIn_1_re; // @[Top.scala 16:14]
  assign fft_io_dIn_1_im = io_dIn_1_im; // @[Top.scala 16:14]
  assign fft_io_din_valid = io_din_valid; // @[Top.scala 17:20]
endmodule
